
module tausworthe_0 ( clock, re_set, tausout );
  output [31:0] tausout;
  input clock, re_set;
  wire   N44, N45, N46, N78, N108, N110, n36, n37, n38, n39, n40, n41, n42,
         n43, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147;
  wire   [31:0] Seed_0;
  wire   [31:0] Seed_1;
  wire   [31:0] Seed_2;
  tri   clock;

  FDS2 \Seed_1_reg[31]  ( .CR(n147), .D(Seed_1[27]), .CP(clock), .QN(n103) );
  FDS2 \Seed_1_reg[28]  ( .CR(n147), .D(Seed_1[24]), .CP(clock), .QN(n106) );
  FDS2 \Seed_1_reg[29]  ( .CR(n147), .D(Seed_1[25]), .CP(clock), .QN(n105) );
  FDS2 \Seed_1_reg[30]  ( .CR(n147), .D(Seed_1[26]), .CP(clock), .QN(n104) );
  FDS2 \Seed_2_reg[21]  ( .CR(n147), .D(Seed_2[4]), .CP(clock), .QN(n89) );
  FDS2 \Seed_2_reg[27]  ( .CR(n147), .D(Seed_2[10]), .CP(clock), .QN(n83) );
  FDS2 \Seed_2_reg[16]  ( .CR(n147), .D(n119), .CP(clock), .QN(n94) );
  FDS2 \Seed_2_reg[22]  ( .CR(n147), .D(Seed_2[5]), .CP(clock), .QN(n88) );
  FDS2 \Seed_2_reg[28]  ( .CR(n147), .D(Seed_2[11]), .CP(clock), .QN(n82) );
  FDS2 \Seed_2_reg[17]  ( .CR(n147), .D(n126), .CP(clock), .QN(n93) );
  FDS2 \Seed_2_reg[23]  ( .CR(n147), .D(Seed_2[6]), .CP(clock), .QN(n87) );
  FDS2 \Seed_2_reg[29]  ( .CR(n147), .D(Seed_2[12]), .CP(clock), .QN(n81) );
  FDS2 \Seed_2_reg[18]  ( .CR(n147), .D(n133), .CP(clock), .QN(n92) );
  FDS2 \Seed_2_reg[24]  ( .CR(n147), .D(Seed_2[7]), .CP(clock), .QN(n86) );
  FDS2 \Seed_2_reg[30]  ( .CR(n147), .D(Seed_2[13]), .CP(clock), .QN(n80) );
  FDS2 \Seed_2_reg[19]  ( .CR(n147), .D(n120), .CP(clock), .QN(n91) );
  FDS2 \Seed_2_reg[25]  ( .CR(n147), .D(Seed_2[8]), .CP(clock), .QN(n85) );
  FDS2 \Seed_2_reg[31]  ( .CR(n147), .D(Seed_2[14]), .CP(clock), .QN(n79) );
  FDS2 \Seed_2_reg[20]  ( .CR(n147), .D(n127), .CP(clock), .QN(n90) );
  FDS2 \Seed_2_reg[26]  ( .CR(n147), .D(Seed_2[9]), .CP(clock), .QN(n84) );
  FDS2 \Seed_2_reg[15]  ( .CR(n147), .D(n131), .CP(clock), .QN(n95) );
  FDS2 \Seed_2_reg[3]  ( .CR(n147), .D(n125), .CP(clock), .QN(n54) );
  FD1 \Seed_2_reg[2]  ( .D(N46), .CP(clock), .QN(n56) );
  FD1 \Seed_2_reg[1]  ( .D(N45), .CP(clock), .QN(n58) );
  FD1 \Seed_2_reg[0]  ( .D(N44), .CP(clock), .QN(n60) );
  FDS2 \Seed_0_reg[25]  ( .CR(n147), .D(Seed_0[13]), .CP(clock), .QN(n67) );
  FDS2 \Seed_0_reg[31]  ( .CR(n147), .D(Seed_0[19]), .CP(clock), .QN(n61) );
  FDS2 \Seed_0_reg[24]  ( .CR(n147), .D(Seed_0[12]), .CP(clock), .QN(n68) );
  FDS2 \Seed_0_reg[30]  ( .CR(n147), .D(Seed_0[18]), .CP(clock), .QN(n62) );
  FDS2 \Seed_0_reg[23]  ( .CR(n147), .D(Seed_0[11]), .CP(clock), .QN(n70) );
  FDS2 \Seed_0_reg[29]  ( .CR(n147), .D(Seed_0[17]), .CP(clock), .QN(n63) );
  FDS2 \Seed_0_reg[22]  ( .CR(n147), .D(Seed_0[10]), .CP(clock), .QN(n73) );
  FDS2 \Seed_0_reg[28]  ( .CR(n147), .D(Seed_0[16]), .CP(clock), .QN(n64) );
  FDS2 \Seed_0_reg[21]  ( .CR(n147), .D(Seed_0[9]), .CP(clock), .QN(n75) );
  FDS2 \Seed_0_reg[27]  ( .CR(n147), .D(Seed_0[15]), .CP(clock), .QN(n65) );
  FDS2 \Seed_0_reg[20]  ( .CR(n147), .D(Seed_0[8]), .CP(clock), .QN(n77) );
  FDS2 \Seed_0_reg[26]  ( .CR(n147), .D(Seed_0[14]), .CP(clock), .QN(n66) );
  FDS2 \Seed_0_reg[0]  ( .CR(n147), .D(n138), .CP(clock), .QN(n59) );
  FDS2 \Seed_1_reg[7]  ( .CR(n147), .D(Seed_1[3]), .CP(clock), .Q(Seed_1[7]), 
        .QN(n47) );
  FDS2 \Seed_1_reg[23]  ( .CR(n147), .D(Seed_1[19]), .CP(clock), .Q(Seed_1[23]), .QN(n111) );
  FDS2 \Seed_1_reg[27]  ( .CR(n147), .D(Seed_1[23]), .CP(clock), .Q(Seed_1[27]), .QN(n107) );
  FDS2 \Seed_1_reg[24]  ( .CR(n147), .D(Seed_1[20]), .CP(clock), .Q(Seed_1[24]), .QN(n109) );
  FDS2 \Seed_1_reg[25]  ( .CR(n147), .D(Seed_1[21]), .CP(clock), .Q(Seed_1[25]), .QN(n110) );
  FDS2 \Seed_1_reg[6]  ( .CR(n147), .D(n113), .CP(clock), .Q(Seed_1[6]), .QN(
        n48) );
  FDS2 \Seed_1_reg[26]  ( .CR(n147), .D(Seed_1[22]), .CP(clock), .Q(Seed_1[26]), .QN(n108) );
  FD1 \Seed_1_reg[2]  ( .D(N110), .CP(clock), .Q(Seed_1[2]) );
  FDS2 \Seed_1_reg[1]  ( .CR(n147), .D(n114), .CP(clock), .Q(Seed_1[1]) );
  FD1 \Seed_1_reg[0]  ( .D(N108), .CP(clock), .Q(Seed_1[0]) );
  FDS2 \Seed_2_reg[4]  ( .CR(n147), .D(n132), .CP(clock), .Q(Seed_2[4]), .QN(
        n52) );
  FDS2 \Seed_2_reg[10]  ( .CR(n147), .D(n117), .CP(clock), .Q(Seed_2[10]), 
        .QN(n98) );
  FDS2 \Seed_2_reg[5]  ( .CR(n147), .D(n121), .CP(clock), .Q(Seed_2[5]), .QN(
        n50) );
  FDS2 \Seed_2_reg[11]  ( .CR(n147), .D(n123), .CP(clock), .Q(Seed_2[11]), 
        .QN(n101) );
  FDS2 \Seed_2_reg[12]  ( .CR(n147), .D(n130), .CP(clock), .Q(Seed_2[12]), 
        .QN(n99) );
  FDS2 \Seed_2_reg[13]  ( .CR(n147), .D(n118), .CP(clock), .Q(Seed_2[13]), 
        .QN(n97) );
  FDS2 \Seed_2_reg[8]  ( .CR(n147), .D(n122), .CP(clock), .Q(Seed_2[8]), .QN(
        n102) );
  FDS2 \Seed_2_reg[14]  ( .CR(n147), .D(n124), .CP(clock), .Q(Seed_2[14]), 
        .QN(n96) );
  FDS2 \Seed_2_reg[9]  ( .CR(n147), .D(n129), .CP(clock), .Q(Seed_2[9]), .QN(
        n100) );
  FDS2 \Seed_0_reg[1]  ( .CR(n147), .D(n137), .CP(clock), .Q(Seed_0[1]), .QN(
        n57) );
  FDS2 \Seed_0_reg[13]  ( .CR(n147), .D(Seed_0[1]), .CP(clock), .Q(Seed_0[13]), 
        .QN(n42) );
  FDS2 \Seed_0_reg[7]  ( .CR(n147), .D(n135), .CP(clock), .Q(Seed_0[7]), .QN(
        n76) );
  FDS2 \Seed_0_reg[19]  ( .CR(n147), .D(Seed_0[7]), .CP(clock), .Q(Seed_0[19]), 
        .QN(n36) );
  FDS2 \Seed_0_reg[12]  ( .CR(n147), .D(n139), .CP(clock), .Q(Seed_0[12]), 
        .QN(n43) );
  FDS2 \Seed_0_reg[6]  ( .CR(n147), .D(n136), .CP(clock), .Q(Seed_0[6]), .QN(
        n78) );
  FDS2 \Seed_0_reg[18]  ( .CR(n147), .D(Seed_0[6]), .CP(clock), .Q(Seed_0[18]), 
        .QN(n37) );
  FDS2 \Seed_0_reg[11]  ( .CR(n147), .D(n141), .CP(clock), .Q(Seed_0[11]), 
        .QN(n69) );
  FDS2 \Seed_0_reg[5]  ( .CR(n147), .D(n140), .CP(clock), .Q(Seed_0[5]), .QN(
        n49) );
  FDS2 \Seed_0_reg[17]  ( .CR(n147), .D(Seed_0[5]), .CP(clock), .Q(Seed_0[17]), 
        .QN(n38) );
  FDS2 \Seed_0_reg[10]  ( .CR(n147), .D(n143), .CP(clock), .Q(Seed_0[10]), 
        .QN(n71) );
  FDS2 \Seed_0_reg[4]  ( .CR(n147), .D(n142), .CP(clock), .Q(Seed_0[4]), .QN(
        n51) );
  FDS2 \Seed_0_reg[16]  ( .CR(n147), .D(Seed_0[4]), .CP(clock), .Q(Seed_0[16]), 
        .QN(n39) );
  FDS2 \Seed_0_reg[9]  ( .CR(n147), .D(n145), .CP(clock), .Q(Seed_0[9]), .QN(
        n72) );
  FDS2 \Seed_0_reg[3]  ( .CR(n147), .D(n144), .CP(clock), .Q(Seed_0[3]), .QN(
        n53) );
  FDS2 \Seed_0_reg[15]  ( .CR(n147), .D(Seed_0[3]), .CP(clock), .Q(Seed_0[15]), 
        .QN(n40) );
  FDS2 \Seed_0_reg[8]  ( .CR(n147), .D(n146), .CP(clock), .Q(Seed_0[8]), .QN(
        n74) );
  FD1 \Seed_0_reg[2]  ( .D(N78), .CP(clock), .Q(Seed_0[2]), .QN(n55) );
  FDS2 \Seed_0_reg[14]  ( .CR(n147), .D(Seed_0[2]), .CP(clock), .Q(Seed_0[14]), 
        .QN(n41) );
  FDS2 \Seed_1_reg[3]  ( .CR(n147), .D(n115), .CP(clock), .Q(Seed_1[3]) );
  FDS2 \Seed_1_reg[11]  ( .CR(n147), .D(Seed_1[7]), .CP(clock), .Q(Seed_1[11])
         );
  FDS2 \Seed_1_reg[15]  ( .CR(n147), .D(Seed_1[11]), .CP(clock), .Q(Seed_1[15]) );
  FDS2 \Seed_1_reg[19]  ( .CR(n147), .D(Seed_1[15]), .CP(clock), .Q(Seed_1[19]) );
  FDS2 \Seed_1_reg[4]  ( .CR(n147), .D(n112), .CP(clock), .Q(Seed_1[4]) );
  FDS2 \Seed_1_reg[8]  ( .CR(n147), .D(Seed_1[4]), .CP(clock), .Q(Seed_1[8])
         );
  FDS2 \Seed_1_reg[12]  ( .CR(n147), .D(Seed_1[8]), .CP(clock), .Q(Seed_1[12])
         );
  FDS2 \Seed_1_reg[16]  ( .CR(n147), .D(Seed_1[12]), .CP(clock), .Q(Seed_1[16]) );
  FDS2 \Seed_1_reg[20]  ( .CR(n147), .D(Seed_1[16]), .CP(clock), .Q(Seed_1[20]) );
  FDS2 \Seed_1_reg[5]  ( .CR(n147), .D(n116), .CP(clock), .Q(Seed_1[5]) );
  FDS2 \Seed_1_reg[9]  ( .CR(n147), .D(Seed_1[5]), .CP(clock), .Q(Seed_1[9])
         );
  FDS2 \Seed_1_reg[13]  ( .CR(n147), .D(Seed_1[9]), .CP(clock), .Q(Seed_1[13])
         );
  FDS2 \Seed_1_reg[17]  ( .CR(n147), .D(Seed_1[13]), .CP(clock), .Q(Seed_1[17]) );
  FDS2 \Seed_1_reg[21]  ( .CR(n147), .D(Seed_1[17]), .CP(clock), .Q(Seed_1[21]) );
  FDS2 \Seed_1_reg[10]  ( .CR(n147), .D(Seed_1[6]), .CP(clock), .Q(Seed_1[10])
         );
  FDS2 \Seed_1_reg[14]  ( .CR(n147), .D(Seed_1[10]), .CP(clock), .Q(Seed_1[14]) );
  FDS2 \Seed_1_reg[18]  ( .CR(n147), .D(Seed_1[14]), .CP(clock), .Q(Seed_1[18]) );
  FDS2 \Seed_1_reg[22]  ( .CR(n147), .D(Seed_1[18]), .CP(clock), .Q(Seed_1[22]) );
  FDS2 \Seed_2_reg[6]  ( .CR(n147), .D(n128), .CP(clock), .Q(Seed_2[6]) );
  FDS2 \Seed_2_reg[7]  ( .CR(n147), .D(n134), .CP(clock), .Q(Seed_2[7]) );
  EO U3 ( .A(n1), .B(n100), .Z(tausout[9]) );
  EO U4 ( .A(Seed_1[9]), .B(n72), .Z(n1) );
  EO U5 ( .A(n2), .B(n102), .Z(tausout[8]) );
  EO U6 ( .A(Seed_1[8]), .B(n74), .Z(n2) );
  EO U7 ( .A(n3), .B(n76), .Z(tausout[7]) );
  EO U8 ( .A(Seed_2[7]), .B(n47), .Z(n3) );
  EO U9 ( .A(n4), .B(n78), .Z(tausout[6]) );
  EO U10 ( .A(Seed_2[6]), .B(n48), .Z(n4) );
  EO U11 ( .A(n5), .B(n50), .Z(tausout[5]) );
  EO U12 ( .A(Seed_1[5]), .B(n49), .Z(n5) );
  EO U13 ( .A(n6), .B(n52), .Z(tausout[4]) );
  EO U14 ( .A(Seed_1[4]), .B(n51), .Z(n6) );
  EO U15 ( .A(n7), .B(n54), .Z(tausout[3]) );
  EO U16 ( .A(Seed_1[3]), .B(n53), .Z(n7) );
  EN U17 ( .A(n103), .B(n8), .Z(tausout[31]) );
  EO U18 ( .A(n61), .B(n79), .Z(n8) );
  EN U19 ( .A(n104), .B(n9), .Z(tausout[30]) );
  EO U20 ( .A(n62), .B(n80), .Z(n9) );
  EO U21 ( .A(n10), .B(n56), .Z(tausout[2]) );
  EO U22 ( .A(Seed_1[2]), .B(n55), .Z(n10) );
  EN U23 ( .A(n105), .B(n11), .Z(tausout[29]) );
  EO U24 ( .A(n63), .B(n81), .Z(n11) );
  EN U25 ( .A(n106), .B(n12), .Z(tausout[28]) );
  EO U26 ( .A(n64), .B(n82), .Z(n12) );
  EN U27 ( .A(n107), .B(n13), .Z(tausout[27]) );
  EO U28 ( .A(n65), .B(n83), .Z(n13) );
  EN U29 ( .A(n108), .B(n14), .Z(tausout[26]) );
  EO U30 ( .A(n66), .B(n84), .Z(n14) );
  EN U31 ( .A(n110), .B(n15), .Z(tausout[25]) );
  EO U32 ( .A(n67), .B(n85), .Z(n15) );
  EN U33 ( .A(n109), .B(n16), .Z(tausout[24]) );
  EO U34 ( .A(n68), .B(n86), .Z(n16) );
  EN U35 ( .A(n111), .B(n17), .Z(tausout[23]) );
  EO U36 ( .A(n70), .B(n87), .Z(n17) );
  EO U37 ( .A(n18), .B(n88), .Z(tausout[22]) );
  EO U38 ( .A(Seed_1[22]), .B(n73), .Z(n18) );
  EO U39 ( .A(n19), .B(n89), .Z(tausout[21]) );
  EO U40 ( .A(Seed_1[21]), .B(n75), .Z(n19) );
  EO U41 ( .A(n20), .B(n90), .Z(tausout[20]) );
  EO U42 ( .A(Seed_1[20]), .B(n77), .Z(n20) );
  EO U43 ( .A(n21), .B(n58), .Z(tausout[1]) );
  EO U44 ( .A(Seed_1[1]), .B(n57), .Z(n21) );
  EO U45 ( .A(n22), .B(n36), .Z(tausout[19]) );
  EO U46 ( .A(Seed_1[19]), .B(n91), .Z(n22) );
  EO U47 ( .A(n23), .B(n37), .Z(tausout[18]) );
  EO U48 ( .A(Seed_1[18]), .B(n92), .Z(n23) );
  EO U49 ( .A(n24), .B(n38), .Z(tausout[17]) );
  EO U50 ( .A(Seed_1[17]), .B(n93), .Z(n24) );
  EO U51 ( .A(n25), .B(n39), .Z(tausout[16]) );
  EO U52 ( .A(Seed_1[16]), .B(n94), .Z(n25) );
  EO U53 ( .A(n26), .B(n40), .Z(tausout[15]) );
  EO U54 ( .A(Seed_1[15]), .B(n95), .Z(n26) );
  EO U55 ( .A(n27), .B(n41), .Z(tausout[14]) );
  EO U56 ( .A(Seed_1[14]), .B(n96), .Z(n27) );
  EO U57 ( .A(n28), .B(n42), .Z(tausout[13]) );
  EO U58 ( .A(Seed_1[13]), .B(n97), .Z(n28) );
  EO U59 ( .A(n29), .B(n43), .Z(tausout[12]) );
  EO U60 ( .A(Seed_1[12]), .B(n99), .Z(n29) );
  EO U61 ( .A(n30), .B(n101), .Z(tausout[11]) );
  EO U62 ( .A(Seed_1[11]), .B(n69), .Z(n30) );
  EO U63 ( .A(n31), .B(n98), .Z(tausout[10]) );
  EO U64 ( .A(Seed_1[10]), .B(n71), .Z(n31) );
  EO U65 ( .A(n32), .B(n60), .Z(tausout[0]) );
  EO U66 ( .A(Seed_1[0]), .B(n59), .Z(n32) );
  EO U67 ( .A(n105), .B(n107), .Z(n112) );
  EO U68 ( .A(n103), .B(n105), .Z(n113) );
  EO U69 ( .A(n108), .B(n109), .Z(n114) );
  EO U70 ( .A(n106), .B(n108), .Z(n115) );
  EO U71 ( .A(n104), .B(n106), .Z(n116) );
  EO U72 ( .A(n89), .B(n92), .Z(n117) );
  EO U73 ( .A(n86), .B(n89), .Z(n118) );
  EO U74 ( .A(n83), .B(n86), .Z(n119) );
  EO U75 ( .A(n80), .B(n83), .Z(n120) );
  EO U76 ( .A(n94), .B(n97), .Z(n121) );
  EO U77 ( .A(n91), .B(n94), .Z(n122) );
  EO U78 ( .A(n88), .B(n91), .Z(n123) );
  EO U79 ( .A(n85), .B(n88), .Z(n124) );
  EO U80 ( .A(n96), .B(n101), .Z(n125) );
  EO U81 ( .A(n82), .B(n85), .Z(n126) );
  EO U82 ( .A(n79), .B(n82), .Z(n127) );
  EO U83 ( .A(n93), .B(n96), .Z(n128) );
  EO U84 ( .A(n90), .B(n93), .Z(n129) );
  EO U85 ( .A(n87), .B(n90), .Z(n130) );
  EO U86 ( .A(n84), .B(n87), .Z(n131) );
  EO U87 ( .A(n95), .B(n99), .Z(n132) );
  EO U88 ( .A(n81), .B(n84), .Z(n133) );
  EO U89 ( .A(n92), .B(n95), .Z(n134) );
  EO U90 ( .A(n66), .B(n42), .Z(n135) );
  EO U91 ( .A(n67), .B(n43), .Z(n136) );
  EO U92 ( .A(n76), .B(n77), .Z(n137) );
  EO U93 ( .A(n78), .B(n36), .Z(n138) );
  EO U94 ( .A(n61), .B(n37), .Z(n139) );
  EO U95 ( .A(n68), .B(n69), .Z(n140) );
  EO U96 ( .A(n62), .B(n38), .Z(n141) );
  EO U97 ( .A(n70), .B(n71), .Z(n142) );
  EO U98 ( .A(n63), .B(n39), .Z(n143) );
  EO U99 ( .A(n72), .B(n73), .Z(n144) );
  EO U100 ( .A(n64), .B(n40), .Z(n145) );
  EO U101 ( .A(n65), .B(n41), .Z(n146) );
  ND2 U102 ( .A(n33), .B(n147), .Z(N78) );
  EN U103 ( .A(n75), .B(n74), .Z(n33) );
  ND2 U104 ( .A(n34), .B(n147), .Z(N46) );
  EN U105 ( .A(n98), .B(n97), .Z(n34) );
  ND2 U106 ( .A(n35), .B(n147), .Z(N45) );
  EN U107 ( .A(n100), .B(n99), .Z(n35) );
  ND2 U108 ( .A(n44), .B(n147), .Z(N44) );
  EN U109 ( .A(n102), .B(n101), .Z(n44) );
  ND2 U110 ( .A(n45), .B(n147), .Z(N110) );
  EN U111 ( .A(n110), .B(n107), .Z(n45) );
  ND2 U112 ( .A(n46), .B(n147), .Z(N108) );
  IV U113 ( .A(re_set), .Z(n147) );
  EN U114 ( .A(n111), .B(n110), .Z(n46) );
endmodule


module tausworthe_1 ( clock, re_set, tausout );
  output [31:0] tausout;
  input clock, re_set;
  wire   N44, N45, N46, N78, N108, N110, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155;
  wire   [31:0] Seed_0;
  wire   [31:0] Seed_1;
  wire   [31:0] Seed_2;
  tri   clock;

  FDS2 \Seed_1_reg[31]  ( .CR(n147), .D(Seed_1[27]), .CP(clock), .QN(n103) );
  FDS2 \Seed_1_reg[28]  ( .CR(n147), .D(Seed_1[24]), .CP(clock), .QN(n106) );
  FDS2 \Seed_1_reg[29]  ( .CR(n147), .D(Seed_1[25]), .CP(clock), .QN(n105) );
  FDS2 \Seed_1_reg[30]  ( .CR(n147), .D(Seed_1[26]), .CP(clock), .QN(n104) );
  FDS2 \Seed_2_reg[21]  ( .CR(n147), .D(Seed_2[4]), .CP(clock), .QN(n89) );
  FDS2 \Seed_2_reg[27]  ( .CR(n147), .D(Seed_2[10]), .CP(clock), .QN(n83) );
  FDS2 \Seed_2_reg[16]  ( .CR(n147), .D(n119), .CP(clock), .QN(n94) );
  FDS2 \Seed_2_reg[22]  ( .CR(n147), .D(Seed_2[5]), .CP(clock), .QN(n88) );
  FDS2 \Seed_2_reg[28]  ( .CR(n147), .D(Seed_2[11]), .CP(clock), .QN(n82) );
  FDS2 \Seed_2_reg[17]  ( .CR(n147), .D(n126), .CP(clock), .QN(n93) );
  FDS2 \Seed_2_reg[23]  ( .CR(n147), .D(Seed_2[6]), .CP(clock), .QN(n87) );
  FDS2 \Seed_2_reg[29]  ( .CR(n147), .D(Seed_2[12]), .CP(clock), .QN(n81) );
  FDS2 \Seed_2_reg[18]  ( .CR(n147), .D(n133), .CP(clock), .QN(n92) );
  FDS2 \Seed_2_reg[24]  ( .CR(n147), .D(Seed_2[7]), .CP(clock), .QN(n86) );
  FDS2 \Seed_2_reg[30]  ( .CR(n147), .D(Seed_2[13]), .CP(clock), .QN(n80) );
  FDS2 \Seed_2_reg[19]  ( .CR(n147), .D(n120), .CP(clock), .QN(n91) );
  FDS2 \Seed_2_reg[25]  ( .CR(n147), .D(Seed_2[8]), .CP(clock), .QN(n85) );
  FDS2 \Seed_2_reg[31]  ( .CR(n147), .D(Seed_2[14]), .CP(clock), .QN(n79) );
  FDS2 \Seed_2_reg[20]  ( .CR(n147), .D(n127), .CP(clock), .QN(n90) );
  FDS2 \Seed_2_reg[26]  ( .CR(n147), .D(Seed_2[9]), .CP(clock), .QN(n84) );
  FDS2 \Seed_2_reg[15]  ( .CR(n147), .D(n131), .CP(clock), .QN(n95) );
  FDS2 \Seed_2_reg[3]  ( .CR(n147), .D(n125), .CP(clock), .QN(n54) );
  FD1 \Seed_2_reg[2]  ( .D(N46), .CP(clock), .QN(n56) );
  FD1 \Seed_2_reg[1]  ( .D(N45), .CP(clock), .QN(n58) );
  FD1 \Seed_2_reg[0]  ( .D(N44), .CP(clock), .QN(n60) );
  FDS2 \Seed_0_reg[25]  ( .CR(n147), .D(Seed_0[13]), .CP(clock), .QN(n67) );
  FDS2 \Seed_0_reg[31]  ( .CR(n147), .D(Seed_0[19]), .CP(clock), .QN(n61) );
  FDS2 \Seed_0_reg[24]  ( .CR(n147), .D(Seed_0[12]), .CP(clock), .QN(n68) );
  FDS2 \Seed_0_reg[30]  ( .CR(n147), .D(Seed_0[18]), .CP(clock), .QN(n62) );
  FDS2 \Seed_0_reg[23]  ( .CR(n147), .D(Seed_0[11]), .CP(clock), .QN(n70) );
  FDS2 \Seed_0_reg[29]  ( .CR(n147), .D(Seed_0[17]), .CP(clock), .QN(n63) );
  FDS2 \Seed_0_reg[22]  ( .CR(n147), .D(Seed_0[10]), .CP(clock), .QN(n73) );
  FDS2 \Seed_0_reg[28]  ( .CR(n147), .D(Seed_0[16]), .CP(clock), .QN(n64) );
  FDS2 \Seed_0_reg[21]  ( .CR(n147), .D(Seed_0[9]), .CP(clock), .QN(n75) );
  FDS2 \Seed_0_reg[27]  ( .CR(n147), .D(Seed_0[15]), .CP(clock), .QN(n65) );
  FDS2 \Seed_0_reg[20]  ( .CR(n147), .D(Seed_0[8]), .CP(clock), .QN(n77) );
  FDS2 \Seed_0_reg[26]  ( .CR(n147), .D(Seed_0[14]), .CP(clock), .QN(n66) );
  FDS2 \Seed_0_reg[0]  ( .CR(n147), .D(n138), .CP(clock), .QN(n59) );
  FDS2 \Seed_1_reg[7]  ( .CR(n147), .D(Seed_1[3]), .CP(clock), .Q(Seed_1[7]), 
        .QN(n47) );
  FDS2 \Seed_1_reg[23]  ( .CR(n147), .D(Seed_1[19]), .CP(clock), .Q(Seed_1[23]), .QN(n111) );
  FDS2 \Seed_1_reg[27]  ( .CR(n147), .D(Seed_1[23]), .CP(clock), .Q(Seed_1[27]), .QN(n107) );
  FDS2 \Seed_1_reg[24]  ( .CR(n147), .D(Seed_1[20]), .CP(clock), .Q(Seed_1[24]), .QN(n109) );
  FDS2 \Seed_1_reg[25]  ( .CR(n147), .D(Seed_1[21]), .CP(clock), .Q(Seed_1[25]), .QN(n110) );
  FDS2 \Seed_1_reg[6]  ( .CR(n147), .D(n113), .CP(clock), .Q(Seed_1[6]), .QN(
        n48) );
  FDS2 \Seed_1_reg[26]  ( .CR(n147), .D(Seed_1[22]), .CP(clock), .Q(Seed_1[26]), .QN(n108) );
  FD1 \Seed_1_reg[2]  ( .D(N110), .CP(clock), .Q(Seed_1[2]) );
  FDS2 \Seed_1_reg[1]  ( .CR(n147), .D(n114), .CP(clock), .Q(Seed_1[1]) );
  FD1 \Seed_1_reg[0]  ( .D(N108), .CP(clock), .Q(Seed_1[0]) );
  FDS2 \Seed_2_reg[4]  ( .CR(n147), .D(n132), .CP(clock), .Q(Seed_2[4]), .QN(
        n52) );
  FDS2 \Seed_2_reg[10]  ( .CR(n147), .D(n117), .CP(clock), .Q(Seed_2[10]), 
        .QN(n98) );
  FDS2 \Seed_2_reg[5]  ( .CR(n147), .D(n121), .CP(clock), .Q(Seed_2[5]), .QN(
        n50) );
  FDS2 \Seed_2_reg[11]  ( .CR(n147), .D(n123), .CP(clock), .Q(Seed_2[11]), 
        .QN(n101) );
  FDS2 \Seed_2_reg[12]  ( .CR(n147), .D(n130), .CP(clock), .Q(Seed_2[12]), 
        .QN(n99) );
  FDS2 \Seed_2_reg[13]  ( .CR(n147), .D(n118), .CP(clock), .Q(Seed_2[13]), 
        .QN(n97) );
  FDS2 \Seed_2_reg[8]  ( .CR(n147), .D(n122), .CP(clock), .Q(Seed_2[8]), .QN(
        n102) );
  FDS2 \Seed_2_reg[14]  ( .CR(n147), .D(n124), .CP(clock), .Q(Seed_2[14]), 
        .QN(n96) );
  FDS2 \Seed_2_reg[9]  ( .CR(n147), .D(n129), .CP(clock), .Q(Seed_2[9]), .QN(
        n100) );
  FDS2 \Seed_0_reg[1]  ( .CR(n147), .D(n137), .CP(clock), .Q(Seed_0[1]), .QN(
        n57) );
  FDS2 \Seed_0_reg[13]  ( .CR(n147), .D(Seed_0[1]), .CP(clock), .Q(Seed_0[13]), 
        .QN(n149) );
  FDS2 \Seed_0_reg[7]  ( .CR(n147), .D(n135), .CP(clock), .Q(Seed_0[7]), .QN(
        n76) );
  FDS2 \Seed_0_reg[19]  ( .CR(n147), .D(Seed_0[7]), .CP(clock), .Q(Seed_0[19]), 
        .QN(n155) );
  FDS2 \Seed_0_reg[12]  ( .CR(n147), .D(n139), .CP(clock), .Q(Seed_0[12]), 
        .QN(n148) );
  FDS2 \Seed_0_reg[6]  ( .CR(n147), .D(n136), .CP(clock), .Q(Seed_0[6]), .QN(
        n78) );
  FDS2 \Seed_0_reg[18]  ( .CR(n147), .D(Seed_0[6]), .CP(clock), .Q(Seed_0[18]), 
        .QN(n154) );
  FDS2 \Seed_0_reg[11]  ( .CR(n147), .D(n141), .CP(clock), .Q(Seed_0[11]), 
        .QN(n69) );
  FDS2 \Seed_0_reg[5]  ( .CR(n147), .D(n140), .CP(clock), .Q(Seed_0[5]), .QN(
        n49) );
  FDS2 \Seed_0_reg[17]  ( .CR(n147), .D(Seed_0[5]), .CP(clock), .Q(Seed_0[17]), 
        .QN(n153) );
  FDS2 \Seed_0_reg[10]  ( .CR(n147), .D(n143), .CP(clock), .Q(Seed_0[10]), 
        .QN(n71) );
  FDS2 \Seed_0_reg[4]  ( .CR(n147), .D(n142), .CP(clock), .Q(Seed_0[4]), .QN(
        n51) );
  FDS2 \Seed_0_reg[16]  ( .CR(n147), .D(Seed_0[4]), .CP(clock), .Q(Seed_0[16]), 
        .QN(n152) );
  FDS2 \Seed_0_reg[9]  ( .CR(n147), .D(n145), .CP(clock), .Q(Seed_0[9]), .QN(
        n72) );
  FDS2 \Seed_0_reg[3]  ( .CR(n147), .D(n144), .CP(clock), .Q(Seed_0[3]), .QN(
        n53) );
  FDS2 \Seed_0_reg[15]  ( .CR(n147), .D(Seed_0[3]), .CP(clock), .Q(Seed_0[15]), 
        .QN(n151) );
  FDS2 \Seed_0_reg[8]  ( .CR(n147), .D(n146), .CP(clock), .Q(Seed_0[8]), .QN(
        n74) );
  FD1 \Seed_0_reg[2]  ( .D(N78), .CP(clock), .Q(Seed_0[2]), .QN(n55) );
  FDS2 \Seed_0_reg[14]  ( .CR(n147), .D(Seed_0[2]), .CP(clock), .Q(Seed_0[14]), 
        .QN(n150) );
  FDS2 \Seed_1_reg[3]  ( .CR(n147), .D(n115), .CP(clock), .Q(Seed_1[3]) );
  FDS2 \Seed_1_reg[11]  ( .CR(n147), .D(Seed_1[7]), .CP(clock), .Q(Seed_1[11])
         );
  FDS2 \Seed_1_reg[15]  ( .CR(n147), .D(Seed_1[11]), .CP(clock), .Q(Seed_1[15]) );
  FDS2 \Seed_1_reg[19]  ( .CR(n147), .D(Seed_1[15]), .CP(clock), .Q(Seed_1[19]) );
  FDS2 \Seed_1_reg[4]  ( .CR(n147), .D(n112), .CP(clock), .Q(Seed_1[4]) );
  FDS2 \Seed_1_reg[8]  ( .CR(n147), .D(Seed_1[4]), .CP(clock), .Q(Seed_1[8])
         );
  FDS2 \Seed_1_reg[12]  ( .CR(n147), .D(Seed_1[8]), .CP(clock), .Q(Seed_1[12])
         );
  FDS2 \Seed_1_reg[16]  ( .CR(n147), .D(Seed_1[12]), .CP(clock), .Q(Seed_1[16]) );
  FDS2 \Seed_1_reg[20]  ( .CR(n147), .D(Seed_1[16]), .CP(clock), .Q(Seed_1[20]) );
  FDS2 \Seed_1_reg[5]  ( .CR(n147), .D(n116), .CP(clock), .Q(Seed_1[5]) );
  FDS2 \Seed_1_reg[9]  ( .CR(n147), .D(Seed_1[5]), .CP(clock), .Q(Seed_1[9])
         );
  FDS2 \Seed_1_reg[13]  ( .CR(n147), .D(Seed_1[9]), .CP(clock), .Q(Seed_1[13])
         );
  FDS2 \Seed_1_reg[17]  ( .CR(n147), .D(Seed_1[13]), .CP(clock), .Q(Seed_1[17]) );
  FDS2 \Seed_1_reg[21]  ( .CR(n147), .D(Seed_1[17]), .CP(clock), .Q(Seed_1[21]) );
  FDS2 \Seed_1_reg[10]  ( .CR(n147), .D(Seed_1[6]), .CP(clock), .Q(Seed_1[10])
         );
  FDS2 \Seed_1_reg[14]  ( .CR(n147), .D(Seed_1[10]), .CP(clock), .Q(Seed_1[14]) );
  FDS2 \Seed_1_reg[18]  ( .CR(n147), .D(Seed_1[14]), .CP(clock), .Q(Seed_1[18]) );
  FDS2 \Seed_1_reg[22]  ( .CR(n147), .D(Seed_1[18]), .CP(clock), .Q(Seed_1[22]) );
  FDS2 \Seed_2_reg[6]  ( .CR(n147), .D(n128), .CP(clock), .Q(Seed_2[6]) );
  FDS2 \Seed_2_reg[7]  ( .CR(n147), .D(n134), .CP(clock), .Q(Seed_2[7]) );
  EO U3 ( .A(n1), .B(n100), .Z(tausout[9]) );
  EO U4 ( .A(Seed_1[9]), .B(n72), .Z(n1) );
  EO U5 ( .A(n2), .B(n102), .Z(tausout[8]) );
  EO U6 ( .A(Seed_1[8]), .B(n74), .Z(n2) );
  EO U7 ( .A(n3), .B(n76), .Z(tausout[7]) );
  EO U8 ( .A(Seed_2[7]), .B(n47), .Z(n3) );
  EO U9 ( .A(n4), .B(n78), .Z(tausout[6]) );
  EO U10 ( .A(Seed_2[6]), .B(n48), .Z(n4) );
  EO U11 ( .A(n5), .B(n50), .Z(tausout[5]) );
  EO U12 ( .A(Seed_1[5]), .B(n49), .Z(n5) );
  EO U13 ( .A(n6), .B(n52), .Z(tausout[4]) );
  EO U14 ( .A(Seed_1[4]), .B(n51), .Z(n6) );
  EO U15 ( .A(n7), .B(n54), .Z(tausout[3]) );
  EO U16 ( .A(Seed_1[3]), .B(n53), .Z(n7) );
  EN U17 ( .A(n103), .B(n8), .Z(tausout[31]) );
  EO U18 ( .A(n61), .B(n79), .Z(n8) );
  EN U19 ( .A(n104), .B(n9), .Z(tausout[30]) );
  EO U20 ( .A(n62), .B(n80), .Z(n9) );
  EO U21 ( .A(n10), .B(n56), .Z(tausout[2]) );
  EO U22 ( .A(Seed_1[2]), .B(n55), .Z(n10) );
  EN U23 ( .A(n105), .B(n11), .Z(tausout[29]) );
  EO U24 ( .A(n63), .B(n81), .Z(n11) );
  EN U25 ( .A(n106), .B(n12), .Z(tausout[28]) );
  EO U26 ( .A(n64), .B(n82), .Z(n12) );
  EN U27 ( .A(n107), .B(n13), .Z(tausout[27]) );
  EO U28 ( .A(n65), .B(n83), .Z(n13) );
  EN U29 ( .A(n108), .B(n14), .Z(tausout[26]) );
  EO U30 ( .A(n66), .B(n84), .Z(n14) );
  EN U31 ( .A(n110), .B(n15), .Z(tausout[25]) );
  EO U32 ( .A(n67), .B(n85), .Z(n15) );
  EN U33 ( .A(n109), .B(n16), .Z(tausout[24]) );
  EO U34 ( .A(n68), .B(n86), .Z(n16) );
  EN U35 ( .A(n111), .B(n17), .Z(tausout[23]) );
  EO U36 ( .A(n70), .B(n87), .Z(n17) );
  EO U37 ( .A(n18), .B(n88), .Z(tausout[22]) );
  EO U38 ( .A(Seed_1[22]), .B(n73), .Z(n18) );
  EO U39 ( .A(n19), .B(n89), .Z(tausout[21]) );
  EO U40 ( .A(Seed_1[21]), .B(n75), .Z(n19) );
  EO U41 ( .A(n20), .B(n90), .Z(tausout[20]) );
  EO U42 ( .A(Seed_1[20]), .B(n77), .Z(n20) );
  EO U43 ( .A(n21), .B(n58), .Z(tausout[1]) );
  EO U44 ( .A(Seed_1[1]), .B(n57), .Z(n21) );
  EO U45 ( .A(n22), .B(n155), .Z(tausout[19]) );
  EO U46 ( .A(Seed_1[19]), .B(n91), .Z(n22) );
  EO U47 ( .A(n23), .B(n154), .Z(tausout[18]) );
  EO U48 ( .A(Seed_1[18]), .B(n92), .Z(n23) );
  EO U49 ( .A(n24), .B(n153), .Z(tausout[17]) );
  EO U50 ( .A(Seed_1[17]), .B(n93), .Z(n24) );
  EO U51 ( .A(n25), .B(n152), .Z(tausout[16]) );
  EO U52 ( .A(Seed_1[16]), .B(n94), .Z(n25) );
  EO U53 ( .A(n26), .B(n151), .Z(tausout[15]) );
  EO U54 ( .A(Seed_1[15]), .B(n95), .Z(n26) );
  EO U55 ( .A(n27), .B(n150), .Z(tausout[14]) );
  EO U56 ( .A(Seed_1[14]), .B(n96), .Z(n27) );
  EO U57 ( .A(n28), .B(n149), .Z(tausout[13]) );
  EO U58 ( .A(Seed_1[13]), .B(n97), .Z(n28) );
  EO U59 ( .A(n29), .B(n148), .Z(tausout[12]) );
  EO U60 ( .A(Seed_1[12]), .B(n99), .Z(n29) );
  EO U61 ( .A(n30), .B(n101), .Z(tausout[11]) );
  EO U62 ( .A(Seed_1[11]), .B(n69), .Z(n30) );
  EO U63 ( .A(n31), .B(n98), .Z(tausout[10]) );
  EO U64 ( .A(Seed_1[10]), .B(n71), .Z(n31) );
  EO U65 ( .A(n32), .B(n60), .Z(tausout[0]) );
  EO U66 ( .A(Seed_1[0]), .B(n59), .Z(n32) );
  EO U67 ( .A(n105), .B(n107), .Z(n112) );
  EO U68 ( .A(n103), .B(n105), .Z(n113) );
  EO U69 ( .A(n108), .B(n109), .Z(n114) );
  EO U70 ( .A(n106), .B(n108), .Z(n115) );
  EO U71 ( .A(n104), .B(n106), .Z(n116) );
  EO U72 ( .A(n89), .B(n92), .Z(n117) );
  EO U73 ( .A(n86), .B(n89), .Z(n118) );
  EO U74 ( .A(n83), .B(n86), .Z(n119) );
  EO U75 ( .A(n80), .B(n83), .Z(n120) );
  EO U76 ( .A(n94), .B(n97), .Z(n121) );
  EO U77 ( .A(n91), .B(n94), .Z(n122) );
  EO U78 ( .A(n88), .B(n91), .Z(n123) );
  EO U79 ( .A(n85), .B(n88), .Z(n124) );
  EO U80 ( .A(n96), .B(n101), .Z(n125) );
  EO U81 ( .A(n82), .B(n85), .Z(n126) );
  EO U82 ( .A(n79), .B(n82), .Z(n127) );
  EO U83 ( .A(n93), .B(n96), .Z(n128) );
  EO U84 ( .A(n90), .B(n93), .Z(n129) );
  EO U85 ( .A(n87), .B(n90), .Z(n130) );
  EO U86 ( .A(n84), .B(n87), .Z(n131) );
  EO U87 ( .A(n95), .B(n99), .Z(n132) );
  EO U88 ( .A(n81), .B(n84), .Z(n133) );
  EO U89 ( .A(n92), .B(n95), .Z(n134) );
  EO U90 ( .A(n66), .B(n149), .Z(n135) );
  EO U91 ( .A(n67), .B(n148), .Z(n136) );
  EO U92 ( .A(n76), .B(n77), .Z(n137) );
  EO U93 ( .A(n78), .B(n155), .Z(n138) );
  EO U94 ( .A(n61), .B(n154), .Z(n139) );
  EO U95 ( .A(n68), .B(n69), .Z(n140) );
  EO U96 ( .A(n62), .B(n153), .Z(n141) );
  EO U97 ( .A(n70), .B(n71), .Z(n142) );
  EO U98 ( .A(n63), .B(n152), .Z(n143) );
  EO U99 ( .A(n72), .B(n73), .Z(n144) );
  EO U100 ( .A(n64), .B(n151), .Z(n145) );
  EO U101 ( .A(n65), .B(n150), .Z(n146) );
  ND2 U102 ( .A(n33), .B(n147), .Z(N78) );
  EN U103 ( .A(n75), .B(n74), .Z(n33) );
  ND2 U104 ( .A(n34), .B(n147), .Z(N46) );
  EN U105 ( .A(n98), .B(n97), .Z(n34) );
  ND2 U106 ( .A(n35), .B(n147), .Z(N45) );
  EN U107 ( .A(n100), .B(n99), .Z(n35) );
  ND2 U108 ( .A(n44), .B(n147), .Z(N44) );
  EN U109 ( .A(n102), .B(n101), .Z(n44) );
  ND2 U110 ( .A(n45), .B(n147), .Z(N110) );
  EN U111 ( .A(n110), .B(n107), .Z(n45) );
  ND2 U112 ( .A(n46), .B(n147), .Z(N108) );
  IV U113 ( .A(re_set), .Z(n147) );
  EN U114 ( .A(n111), .B(n110), .Z(n46) );
endmodule


module Poly_Logarithm_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [24:0] carry;
  assign DIFF[0] = B[0];

  FA1A U2_21 ( .A(A[21]), .B(n3), .CI(carry[21]), .CO(carry[22]), .S(DIFF[21])
         );
  FA1A U2_20 ( .A(A[20]), .B(n4), .CI(carry[20]), .CO(carry[21]), .S(DIFF[20])
         );
  FA1A U2_19 ( .A(A[19]), .B(n5), .CI(carry[19]), .CO(carry[20]), .S(DIFF[19])
         );
  FA1A U2_18 ( .A(A[18]), .B(n6), .CI(carry[18]), .CO(carry[19]), .S(DIFF[18])
         );
  FA1A U2_17 ( .A(A[17]), .B(n7), .CI(carry[17]), .CO(carry[18]), .S(DIFF[17])
         );
  FA1A U2_16 ( .A(A[16]), .B(n8), .CI(carry[16]), .CO(carry[17]), .S(DIFF[16])
         );
  FA1A U2_15 ( .A(A[15]), .B(n9), .CI(carry[15]), .CO(carry[16]), .S(DIFF[15])
         );
  FA1A U2_14 ( .A(A[14]), .B(n10), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  FA1A U2_13 ( .A(A[13]), .B(n11), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  FA1A U2_22 ( .A(A[22]), .B(n2), .CI(carry[22]), .CO(carry[23]), .S(DIFF[22])
         );
  EO U1 ( .A(n23), .B(n24), .Z(DIFF[1]) );
  EO U2 ( .A(n22), .B(carry[2]), .Z(DIFF[2]) );
  EO U3 ( .A(n21), .B(carry[3]), .Z(DIFF[3]) );
  EO U4 ( .A(n20), .B(carry[4]), .Z(DIFF[4]) );
  EO U5 ( .A(n19), .B(carry[5]), .Z(DIFF[5]) );
  EO U6 ( .A(n18), .B(carry[6]), .Z(DIFF[6]) );
  EO U7 ( .A(n17), .B(carry[7]), .Z(DIFF[7]) );
  EO U8 ( .A(n16), .B(carry[8]), .Z(DIFF[8]) );
  EO U9 ( .A(n15), .B(carry[9]), .Z(DIFF[9]) );
  EO U10 ( .A(n14), .B(carry[10]), .Z(DIFF[10]) );
  EO U11 ( .A(n13), .B(carry[11]), .Z(DIFF[11]) );
  EO U12 ( .A(n12), .B(carry[12]), .Z(DIFF[12]) );
  IVP U13 ( .A(carry[23]), .Z(DIFF[23]) );
  IVP U14 ( .A(B[22]), .Z(n2) );
  IVP U15 ( .A(B[13]), .Z(n11) );
  IVP U16 ( .A(B[14]), .Z(n10) );
  IVP U17 ( .A(B[15]), .Z(n9) );
  IVP U18 ( .A(B[16]), .Z(n8) );
  IVP U19 ( .A(B[17]), .Z(n7) );
  IVP U20 ( .A(B[18]), .Z(n6) );
  IVP U21 ( .A(B[19]), .Z(n5) );
  IVP U22 ( .A(B[20]), .Z(n4) );
  IVP U23 ( .A(B[21]), .Z(n3) );
  IVP U24 ( .A(B[0]), .Z(n24) );
  IVP U25 ( .A(B[1]), .Z(n23) );
  IVP U26 ( .A(B[2]), .Z(n22) );
  IVP U27 ( .A(B[3]), .Z(n21) );
  IVP U28 ( .A(B[4]), .Z(n20) );
  IVP U29 ( .A(B[5]), .Z(n19) );
  IVP U30 ( .A(B[6]), .Z(n18) );
  IVP U31 ( .A(B[7]), .Z(n17) );
  IVP U32 ( .A(B[8]), .Z(n16) );
  IVP U33 ( .A(B[9]), .Z(n15) );
  IVP U34 ( .A(B[10]), .Z(n14) );
  IVP U35 ( .A(B[11]), .Z(n13) );
  IVP U36 ( .A(B[12]), .Z(n12) );
  AN2P U37 ( .A(n14), .B(carry[10]), .Z(carry[11]) );
  AN2P U38 ( .A(n13), .B(carry[11]), .Z(carry[12]) );
  AN2P U39 ( .A(n12), .B(carry[12]), .Z(carry[13]) );
  AN2P U40 ( .A(n23), .B(n24), .Z(carry[2]) );
  AN2P U41 ( .A(n22), .B(carry[2]), .Z(carry[3]) );
  AN2P U42 ( .A(n21), .B(carry[3]), .Z(carry[4]) );
  AN2P U43 ( .A(n20), .B(carry[4]), .Z(carry[5]) );
  AN2P U44 ( .A(n19), .B(carry[5]), .Z(carry[6]) );
  AN2P U45 ( .A(n18), .B(carry[6]), .Z(carry[7]) );
  AN2P U46 ( .A(n17), .B(carry[7]), .Z(carry[8]) );
  AN2P U47 ( .A(n16), .B(carry[8]), .Z(carry[9]) );
  AN2P U48 ( .A(n15), .B(carry[9]), .Z(carry[10]) );
endmodule


module Poly_Logarithm_DW01_add_2 ( A, B, CI, SUM, CO );
  input [67:0] A;
  input [67:0] B;
  output [67:0] SUM;
  input CI;
  output CO;
  wire   \A[45] , \A[44] , \A[43] , \A[42] , \A[41] , \A[40] , \A[37] , n1, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115;
  assign SUM[46] = A[46];
  assign SUM[39] = A[39];
  assign SUM[38] = A[38];
  assign SUM[36] = A[36];
  assign SUM[45] = \A[45] ;
  assign \A[45]  = A[45];
  assign SUM[44] = \A[44] ;
  assign \A[44]  = A[44];
  assign SUM[43] = \A[43] ;
  assign \A[43]  = A[43];
  assign SUM[42] = \A[42] ;
  assign \A[42]  = A[42];
  assign SUM[41] = \A[41] ;
  assign \A[41]  = A[41];
  assign SUM[40] = \A[40] ;
  assign \A[40]  = A[40];
  assign SUM[37] = \A[37] ;
  assign \A[37]  = A[37];

  OR2P U2 ( .A(B[47]), .B(A[47]), .Z(n1) );
  AN2P U3 ( .A(n1), .B(n115), .Z(SUM[47]) );
  IVP U4 ( .A(n49), .Z(n14) );
  IVP U5 ( .A(n46), .Z(n20) );
  IVP U6 ( .A(n105), .Z(n24) );
  IVP U7 ( .A(n68), .Z(n12) );
  IVP U8 ( .A(n100), .Z(n23) );
  IVP U9 ( .A(n38), .Z(n7) );
  IVP U10 ( .A(n33), .Z(n5) );
  IVP U11 ( .A(n29), .Z(n3) );
  IVP U12 ( .A(n115), .Z(n26) );
  IVP U13 ( .A(n75), .Z(n11) );
  IVP U14 ( .A(n91), .Z(n16) );
  IVP U15 ( .A(n32), .Z(n4) );
  IVP U16 ( .A(n110), .Z(n22) );
  IVP U17 ( .A(n101), .Z(n21) );
  IVP U18 ( .A(n95), .Z(n18) );
  IVP U19 ( .A(n85), .Z(n17) );
  IVP U20 ( .A(n80), .Z(n15) );
  IVP U21 ( .A(n77), .Z(n13) );
  IVP U22 ( .A(n65), .Z(n10) );
  IVP U23 ( .A(n69), .Z(n9) );
  IVP U24 ( .A(n59), .Z(n8) );
  IVP U25 ( .A(n99), .Z(n25) );
  IVP U26 ( .A(n86), .Z(n19) );
  IVP U27 ( .A(n54), .Z(n6) );
  EO U28 ( .A(n27), .B(n28), .Z(SUM[65]) );
  EO U29 ( .A(B[65]), .B(A[65]), .Z(n28) );
  AO7 U30 ( .A(n29), .B(n4), .C(n30), .Z(n27) );
  EO U31 ( .A(n31), .B(n4), .Z(SUM[64]) );
  AO7 U32 ( .A(n33), .B(n34), .C(n35), .Z(n32) );
  AO6 U33 ( .A(n36), .B(n6), .C(n37), .Z(n34) );
  AO7 U34 ( .A(n38), .B(n39), .C(n40), .Z(n36) );
  AO6 U35 ( .A(n41), .B(n8), .C(n42), .Z(n39) );
  AO7 U36 ( .A(n43), .B(n44), .C(n45), .Z(n41) );
  AO1 U37 ( .A(n14), .B(n46), .C(n47), .D(n48), .Z(n43) );
  NR2 U38 ( .A(n49), .B(n50), .Z(n48) );
  ND2 U39 ( .A(n3), .B(n30), .Z(n31) );
  ND2 U40 ( .A(B[64]), .B(A[64]), .Z(n30) );
  NR2 U41 ( .A(B[64]), .B(A[64]), .Z(n29) );
  EO U42 ( .A(n51), .B(n52), .Z(SUM[63]) );
  AO6 U43 ( .A(n53), .B(n6), .C(n37), .Z(n52) );
  ND2 U44 ( .A(n5), .B(n35), .Z(n51) );
  ND2 U45 ( .A(B[63]), .B(A[63]), .Z(n35) );
  NR2 U46 ( .A(B[63]), .B(A[63]), .Z(n33) );
  EO U47 ( .A(n53), .B(n55), .Z(SUM[62]) );
  NR2 U48 ( .A(n37), .B(n54), .Z(n55) );
  NR2 U49 ( .A(B[62]), .B(A[62]), .Z(n54) );
  AN2 U50 ( .A(B[62]), .B(A[62]), .Z(n37) );
  AO7 U51 ( .A(n38), .B(n56), .C(n40), .Z(n53) );
  EO U52 ( .A(n57), .B(n56), .Z(SUM[61]) );
  AO6 U53 ( .A(n8), .B(n58), .C(n42), .Z(n56) );
  ND2 U54 ( .A(n7), .B(n40), .Z(n57) );
  ND2 U55 ( .A(B[61]), .B(A[61]), .Z(n40) );
  NR2 U56 ( .A(B[61]), .B(A[61]), .Z(n38) );
  EO U57 ( .A(n58), .B(n60), .Z(SUM[60]) );
  NR2 U58 ( .A(n42), .B(n59), .Z(n60) );
  NR2 U59 ( .A(B[60]), .B(A[60]), .Z(n59) );
  AN2 U60 ( .A(B[60]), .B(A[60]), .Z(n42) );
  AO7 U61 ( .A(n61), .B(n44), .C(n45), .Z(n58) );
  AO6 U62 ( .A(n9), .B(n62), .C(n63), .Z(n45) );
  AO7 U63 ( .A(n64), .B(n65), .C(n66), .Z(n62) );
  AO6 U64 ( .A(n11), .B(n12), .C(n67), .Z(n64) );
  ND4 U65 ( .A(n9), .B(n10), .C(n11), .D(n13), .Z(n44) );
  EO U66 ( .A(n70), .B(n71), .Z(SUM[59]) );
  NR2 U67 ( .A(n63), .B(n69), .Z(n71) );
  NR2 U68 ( .A(B[59]), .B(A[59]), .Z(n69) );
  AN2 U69 ( .A(B[59]), .B(A[59]), .Z(n63) );
  AO7 U70 ( .A(n65), .B(n72), .C(n66), .Z(n70) );
  EO U71 ( .A(n73), .B(n72), .Z(SUM[58]) );
  AO6 U72 ( .A(n11), .B(n74), .C(n67), .Z(n72) );
  ND2 U73 ( .A(n10), .B(n66), .Z(n73) );
  ND2 U74 ( .A(B[58]), .B(A[58]), .Z(n66) );
  NR2 U75 ( .A(B[58]), .B(A[58]), .Z(n65) );
  EO U76 ( .A(n74), .B(n76), .Z(SUM[57]) );
  NR2 U77 ( .A(n67), .B(n75), .Z(n76) );
  NR2 U78 ( .A(B[57]), .B(A[57]), .Z(n75) );
  AN2 U79 ( .A(B[57]), .B(A[57]), .Z(n67) );
  AO7 U80 ( .A(n77), .B(n61), .C(n68), .Z(n74) );
  EO U81 ( .A(n78), .B(n61), .Z(SUM[56]) );
  AO6 U82 ( .A(n79), .B(n14), .C(n47), .Z(n61) );
  AO7 U83 ( .A(n80), .B(n81), .C(n82), .Z(n47) );
  AO6 U84 ( .A(n83), .B(n16), .C(n84), .Z(n81) );
  AO7 U85 ( .A(n85), .B(n86), .C(n87), .Z(n83) );
  ND4 U86 ( .A(n15), .B(n16), .C(n17), .D(n18), .Z(n49) );
  ND2 U87 ( .A(n13), .B(n68), .Z(n78) );
  ND2 U88 ( .A(B[56]), .B(A[56]), .Z(n68) );
  NR2 U89 ( .A(B[56]), .B(A[56]), .Z(n77) );
  EO U90 ( .A(n88), .B(n89), .Z(SUM[55]) );
  AO6 U91 ( .A(n90), .B(n16), .C(n84), .Z(n89) );
  ND2 U92 ( .A(n15), .B(n82), .Z(n88) );
  ND2 U93 ( .A(B[55]), .B(A[55]), .Z(n82) );
  NR2 U94 ( .A(B[55]), .B(A[55]), .Z(n80) );
  EO U95 ( .A(n90), .B(n92), .Z(SUM[54]) );
  NR2 U96 ( .A(n84), .B(n91), .Z(n92) );
  NR2 U97 ( .A(B[54]), .B(A[54]), .Z(n91) );
  AN2 U98 ( .A(B[54]), .B(A[54]), .Z(n84) );
  AO7 U99 ( .A(n85), .B(n93), .C(n87), .Z(n90) );
  EO U100 ( .A(n94), .B(n93), .Z(SUM[53]) );
  AO6 U101 ( .A(n18), .B(n79), .C(n19), .Z(n93) );
  ND2 U102 ( .A(n17), .B(n87), .Z(n94) );
  ND2 U103 ( .A(B[53]), .B(A[53]), .Z(n87) );
  NR2 U104 ( .A(B[53]), .B(A[53]), .Z(n85) );
  EO U105 ( .A(n79), .B(n96), .Z(SUM[52]) );
  NR2 U106 ( .A(n19), .B(n95), .Z(n96) );
  NR2 U107 ( .A(B[52]), .B(A[52]), .Z(n95) );
  ND2 U108 ( .A(B[52]), .B(A[52]), .Z(n86) );
  ND2 U109 ( .A(n20), .B(n50), .Z(n79) );
  ND4 U110 ( .A(n26), .B(n21), .C(n97), .D(n98), .Z(n50) );
  NR2 U111 ( .A(n99), .B(n100), .Z(n97) );
  AO7 U112 ( .A(n101), .B(n102), .C(n103), .Z(n46) );
  AO6 U113 ( .A(n104), .B(n98), .C(n22), .Z(n102) );
  AO7 U114 ( .A(n100), .B(n105), .C(n106), .Z(n104) );
  EO U115 ( .A(n107), .B(n108), .Z(SUM[51]) );
  AO6 U116 ( .A(n109), .B(n98), .C(n22), .Z(n108) );
  ND2 U117 ( .A(n21), .B(n103), .Z(n107) );
  ND2 U118 ( .A(B[51]), .B(A[51]), .Z(n103) );
  NR2 U119 ( .A(B[51]), .B(A[51]), .Z(n101) );
  EN U120 ( .A(n111), .B(n109), .Z(SUM[50]) );
  AO7 U121 ( .A(n100), .B(n112), .C(n106), .Z(n109) );
  ND2 U122 ( .A(n98), .B(n110), .Z(n111) );
  ND2 U123 ( .A(B[50]), .B(A[50]), .Z(n110) );
  OR2 U124 ( .A(B[50]), .B(A[50]), .Z(n98) );
  EO U125 ( .A(n113), .B(n112), .Z(SUM[49]) );
  AO6 U126 ( .A(n25), .B(n26), .C(n24), .Z(n112) );
  ND2 U127 ( .A(n23), .B(n106), .Z(n113) );
  ND2 U128 ( .A(B[49]), .B(A[49]), .Z(n106) );
  NR2 U129 ( .A(B[49]), .B(A[49]), .Z(n100) );
  EN U130 ( .A(n114), .B(n26), .Z(SUM[48]) );
  ND2 U131 ( .A(n25), .B(n105), .Z(n114) );
  ND2 U132 ( .A(B[48]), .B(A[48]), .Z(n105) );
  NR2 U133 ( .A(B[48]), .B(A[48]), .Z(n99) );
  ND2 U134 ( .A(B[47]), .B(A[47]), .Z(n115) );
endmodule


module Poly_Logarithm_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [47:0] A;
  input [21:0] B;
  output [69:0] PRODUCT;
  input TC;
  wire   \ab[47][21] , \ab[47][20] , \ab[47][19] , \ab[47][18] , \ab[47][17] ,
         \ab[47][16] , \ab[47][15] , \ab[47][14] , \ab[47][13] , \ab[47][12] ,
         \ab[47][11] , \ab[47][10] , \ab[47][9] , \ab[47][8] , \ab[47][7] ,
         \ab[47][6] , \ab[47][5] , \ab[47][4] , \ab[47][3] , \ab[47][2] ,
         \ab[47][1] , \ab[47][0] , \ab[46][21] , \ab[46][20] , \ab[46][19] ,
         \ab[46][18] , \ab[46][17] , \ab[46][16] , \ab[46][15] , \ab[46][14] ,
         \ab[46][13] , \ab[46][12] , \ab[46][11] , \ab[46][10] , \ab[46][9] ,
         \ab[46][8] , \ab[46][7] , \ab[46][6] , \ab[46][5] , \ab[46][4] ,
         \ab[46][3] , \ab[46][2] , \ab[46][1] , \ab[46][0] , \ab[45][21] ,
         \ab[45][20] , \ab[45][19] , \ab[45][18] , \ab[45][17] , \ab[45][16] ,
         \ab[45][15] , \ab[45][14] , \ab[45][13] , \ab[45][12] , \ab[45][11] ,
         \ab[45][10] , \ab[45][9] , \ab[45][8] , \ab[45][7] , \ab[45][6] ,
         \ab[45][5] , \ab[45][4] , \ab[45][3] , \ab[45][2] , \ab[45][1] ,
         \ab[45][0] , \ab[44][21] , \ab[44][20] , \ab[44][19] , \ab[44][18] ,
         \ab[44][17] , \ab[44][16] , \ab[44][15] , \ab[44][14] , \ab[44][13] ,
         \ab[44][12] , \ab[44][11] , \ab[44][10] , \ab[44][9] , \ab[44][8] ,
         \ab[44][7] , \ab[44][6] , \ab[44][5] , \ab[44][4] , \ab[44][3] ,
         \ab[44][2] , \ab[44][1] , \ab[44][0] , \ab[43][21] , \ab[43][20] ,
         \ab[43][19] , \ab[43][18] , \ab[43][17] , \ab[43][16] , \ab[43][15] ,
         \ab[43][14] , \ab[43][13] , \ab[43][12] , \ab[43][11] , \ab[43][10] ,
         \ab[43][9] , \ab[43][8] , \ab[43][7] , \ab[43][6] , \ab[43][5] ,
         \ab[43][4] , \ab[43][3] , \ab[43][2] , \ab[43][1] , \ab[43][0] ,
         \ab[42][21] , \ab[42][20] , \ab[42][19] , \ab[42][18] , \ab[42][17] ,
         \ab[42][16] , \ab[42][15] , \ab[42][14] , \ab[42][13] , \ab[42][12] ,
         \ab[42][11] , \ab[42][10] , \ab[42][9] , \ab[42][8] , \ab[42][7] ,
         \ab[42][6] , \ab[42][5] , \ab[42][4] , \ab[42][3] , \ab[42][2] ,
         \ab[42][1] , \ab[42][0] , \ab[41][21] , \ab[41][20] , \ab[41][19] ,
         \ab[41][18] , \ab[41][17] , \ab[41][16] , \ab[41][15] , \ab[41][14] ,
         \ab[41][13] , \ab[41][12] , \ab[41][11] , \ab[41][10] , \ab[41][9] ,
         \ab[41][8] , \ab[41][7] , \ab[41][6] , \ab[41][5] , \ab[41][4] ,
         \ab[41][3] , \ab[41][2] , \ab[41][1] , \ab[41][0] , \ab[40][21] ,
         \ab[40][20] , \ab[40][19] , \ab[40][18] , \ab[40][17] , \ab[40][16] ,
         \ab[40][15] , \ab[40][14] , \ab[40][13] , \ab[40][12] , \ab[40][11] ,
         \ab[40][10] , \ab[40][9] , \ab[40][8] , \ab[40][7] , \ab[40][6] ,
         \ab[40][5] , \ab[40][4] , \ab[40][3] , \ab[40][2] , \ab[40][1] ,
         \ab[40][0] , \ab[39][21] , \ab[39][20] , \ab[39][19] , \ab[39][18] ,
         \ab[39][17] , \ab[39][16] , \ab[39][15] , \ab[39][14] , \ab[39][13] ,
         \ab[39][12] , \ab[39][11] , \ab[39][10] , \ab[39][9] , \ab[39][8] ,
         \ab[39][7] , \ab[39][6] , \ab[39][5] , \ab[39][4] , \ab[39][3] ,
         \ab[39][2] , \ab[39][1] , \ab[39][0] , \ab[38][21] , \ab[38][20] ,
         \ab[38][19] , \ab[38][18] , \ab[38][17] , \ab[38][16] , \ab[38][15] ,
         \ab[38][14] , \ab[38][13] , \ab[38][12] , \ab[38][11] , \ab[38][10] ,
         \ab[38][9] , \ab[38][8] , \ab[38][7] , \ab[38][6] , \ab[38][5] ,
         \ab[38][4] , \ab[38][3] , \ab[38][2] , \ab[38][1] , \ab[38][0] ,
         \ab[37][21] , \ab[37][20] , \ab[37][19] , \ab[37][18] , \ab[37][17] ,
         \ab[37][16] , \ab[37][15] , \ab[37][14] , \ab[37][13] , \ab[37][12] ,
         \ab[37][11] , \ab[37][10] , \ab[37][9] , \ab[37][8] , \ab[37][7] ,
         \ab[37][6] , \ab[37][5] , \ab[37][4] , \ab[37][3] , \ab[37][2] ,
         \ab[37][1] , \ab[37][0] , \ab[36][21] , \ab[36][20] , \ab[36][19] ,
         \ab[36][18] , \ab[36][17] , \ab[36][16] , \ab[36][15] , \ab[36][14] ,
         \ab[36][13] , \ab[36][12] , \ab[36][11] , \ab[36][10] , \ab[36][9] ,
         \ab[36][8] , \ab[36][7] , \ab[36][6] , \ab[36][5] , \ab[36][4] ,
         \ab[36][3] , \ab[36][2] , \ab[36][1] , \ab[36][0] , \ab[35][21] ,
         \ab[35][20] , \ab[35][19] , \ab[35][18] , \ab[35][17] , \ab[35][16] ,
         \ab[35][15] , \ab[35][14] , \ab[35][13] , \ab[35][12] , \ab[35][11] ,
         \ab[35][10] , \ab[35][9] , \ab[35][8] , \ab[35][7] , \ab[35][6] ,
         \ab[35][5] , \ab[35][4] , \ab[35][3] , \ab[35][2] , \ab[35][1] ,
         \ab[35][0] , \ab[34][21] , \ab[34][20] , \ab[34][19] , \ab[34][18] ,
         \ab[34][17] , \ab[34][16] , \ab[34][15] , \ab[34][14] , \ab[34][13] ,
         \ab[34][12] , \ab[34][11] , \ab[34][10] , \ab[34][9] , \ab[34][8] ,
         \ab[34][7] , \ab[34][6] , \ab[34][5] , \ab[34][4] , \ab[34][3] ,
         \ab[34][2] , \ab[34][1] , \ab[34][0] , \ab[33][21] , \ab[33][20] ,
         \ab[33][19] , \ab[33][18] , \ab[33][17] , \ab[33][16] , \ab[33][15] ,
         \ab[33][14] , \ab[33][13] , \ab[33][12] , \ab[33][11] , \ab[33][10] ,
         \ab[33][9] , \ab[33][8] , \ab[33][7] , \ab[33][6] , \ab[33][5] ,
         \ab[33][4] , \ab[33][3] , \ab[33][2] , \ab[33][1] , \ab[33][0] ,
         \ab[32][21] , \ab[32][20] , \ab[32][19] , \ab[32][18] , \ab[32][17] ,
         \ab[32][16] , \ab[32][15] , \ab[32][14] , \ab[32][13] , \ab[32][12] ,
         \ab[32][11] , \ab[32][10] , \ab[32][9] , \ab[32][8] , \ab[32][7] ,
         \ab[32][6] , \ab[32][5] , \ab[32][4] , \ab[32][3] , \ab[32][2] ,
         \ab[32][1] , \ab[32][0] , \ab[31][21] , \ab[31][20] , \ab[31][19] ,
         \ab[31][18] , \ab[31][17] , \ab[31][16] , \ab[31][15] , \ab[31][14] ,
         \ab[31][13] , \ab[31][12] , \ab[31][11] , \ab[31][10] , \ab[31][9] ,
         \ab[31][8] , \ab[31][7] , \ab[31][6] , \ab[31][5] , \ab[31][4] ,
         \ab[31][3] , \ab[31][2] , \ab[31][1] , \ab[31][0] , \ab[30][21] ,
         \ab[30][20] , \ab[30][19] , \ab[30][18] , \ab[30][17] , \ab[30][16] ,
         \ab[30][15] , \ab[30][14] , \ab[30][13] , \ab[30][12] , \ab[30][11] ,
         \ab[30][10] , \ab[30][9] , \ab[30][8] , \ab[30][7] , \ab[30][6] ,
         \ab[30][5] , \ab[30][4] , \ab[30][3] , \ab[30][2] , \ab[30][1] ,
         \ab[30][0] , \ab[29][21] , \ab[29][20] , \ab[29][19] , \ab[29][18] ,
         \ab[29][17] , \ab[29][16] , \ab[29][15] , \ab[29][14] , \ab[29][13] ,
         \ab[29][12] , \ab[29][11] , \ab[29][10] , \ab[29][9] , \ab[29][8] ,
         \ab[29][7] , \ab[29][6] , \ab[29][5] , \ab[29][4] , \ab[29][3] ,
         \ab[29][2] , \ab[29][1] , \ab[29][0] , \ab[28][21] , \ab[28][20] ,
         \ab[28][19] , \ab[28][18] , \ab[28][17] , \ab[28][16] , \ab[28][15] ,
         \ab[28][14] , \ab[28][13] , \ab[28][12] , \ab[28][11] , \ab[28][10] ,
         \ab[28][9] , \ab[28][8] , \ab[28][7] , \ab[28][6] , \ab[28][5] ,
         \ab[28][4] , \ab[28][3] , \ab[28][2] , \ab[28][1] , \ab[28][0] ,
         \ab[27][21] , \ab[27][20] , \ab[27][19] , \ab[27][18] , \ab[27][17] ,
         \ab[27][16] , \ab[27][15] , \ab[27][14] , \ab[27][13] , \ab[27][12] ,
         \ab[27][11] , \ab[27][10] , \ab[27][9] , \ab[27][8] , \ab[27][7] ,
         \ab[27][6] , \ab[27][5] , \ab[27][4] , \ab[27][3] , \ab[27][2] ,
         \ab[27][1] , \ab[27][0] , \ab[26][21] , \ab[26][20] , \ab[26][19] ,
         \ab[26][18] , \ab[26][17] , \ab[26][16] , \ab[26][15] , \ab[26][14] ,
         \ab[26][13] , \ab[26][12] , \ab[26][11] , \ab[26][10] , \ab[26][9] ,
         \ab[26][8] , \ab[26][7] , \ab[26][6] , \ab[26][5] , \ab[26][4] ,
         \ab[26][3] , \ab[26][2] , \ab[26][1] , \ab[26][0] , \ab[25][21] ,
         \ab[25][20] , \ab[25][19] , \ab[25][18] , \ab[25][17] , \ab[25][16] ,
         \ab[25][15] , \ab[25][14] , \ab[25][13] , \ab[25][12] , \ab[25][11] ,
         \ab[25][10] , \ab[25][9] , \ab[25][8] , \ab[25][7] , \ab[25][6] ,
         \ab[25][5] , \ab[25][4] , \ab[25][3] , \ab[25][2] , \ab[25][1] ,
         \ab[25][0] , \ab[24][21] , \ab[24][20] , \ab[24][19] , \ab[24][18] ,
         \ab[24][17] , \ab[24][16] , \ab[24][15] , \ab[24][14] , \ab[24][13] ,
         \ab[24][12] , \ab[24][11] , \ab[24][10] , \ab[24][9] , \ab[24][8] ,
         \ab[24][7] , \ab[24][6] , \ab[24][5] , \ab[24][4] , \ab[24][3] ,
         \ab[24][2] , \ab[24][1] , \ab[24][0] , \ab[23][21] , \ab[23][20] ,
         \ab[23][19] , \ab[23][18] , \ab[23][17] , \ab[23][16] , \ab[23][15] ,
         \ab[23][14] , \ab[23][13] , \ab[23][12] , \ab[23][11] , \ab[23][10] ,
         \ab[23][9] , \ab[23][8] , \ab[23][7] , \ab[23][6] , \ab[23][5] ,
         \ab[23][4] , \ab[23][3] , \ab[23][2] , \ab[23][1] , \ab[23][0] ,
         \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] , \ab[22][17] ,
         \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] , \ab[22][12] ,
         \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] , \ab[22][7] ,
         \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] , \ab[22][2] ,
         \ab[22][1] , \ab[22][0] , \ab[21][21] , \ab[21][20] , \ab[21][19] ,
         \ab[21][18] , \ab[21][17] , \ab[21][16] , \ab[21][15] , \ab[21][14] ,
         \ab[21][13] , \ab[21][12] , \ab[21][11] , \ab[21][10] , \ab[21][9] ,
         \ab[21][8] , \ab[21][7] , \ab[21][6] , \ab[21][5] , \ab[21][4] ,
         \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][21] ,
         \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] ,
         \ab[20][15] , \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] ,
         \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] ,
         \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] ,
         \ab[20][0] , \ab[19][21] , \ab[19][20] , \ab[19][19] , \ab[19][18] ,
         \ab[19][17] , \ab[19][16] , \ab[19][15] , \ab[19][14] , \ab[19][13] ,
         \ab[19][12] , \ab[19][11] , \ab[19][10] , \ab[19][9] , \ab[19][8] ,
         \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] , \ab[19][3] ,
         \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][21] , \ab[18][20] ,
         \ab[18][19] , \ab[18][18] , \ab[18][17] , \ab[18][16] , \ab[18][15] ,
         \ab[18][14] , \ab[18][13] , \ab[18][12] , \ab[18][11] , \ab[18][10] ,
         \ab[18][9] , \ab[18][8] , \ab[18][7] , \ab[18][6] , \ab[18][5] ,
         \ab[18][4] , \ab[18][3] , \ab[18][2] , \ab[18][1] , \ab[18][0] ,
         \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] , \ab[17][17] ,
         \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] , \ab[17][12] ,
         \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] , \ab[17][7] ,
         \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] , \ab[17][2] ,
         \ab[17][1] , \ab[17][0] , \ab[16][21] , \ab[16][20] , \ab[16][19] ,
         \ab[16][18] , \ab[16][17] , \ab[16][16] , \ab[16][15] , \ab[16][14] ,
         \ab[16][13] , \ab[16][12] , \ab[16][11] , \ab[16][10] , \ab[16][9] ,
         \ab[16][8] , \ab[16][7] , \ab[16][6] , \ab[16][5] , \ab[16][4] ,
         \ab[16][3] , \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][21] ,
         \ab[15][20] , \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] ,
         \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][21] , \ab[14][20] , \ab[14][19] , \ab[14][18] ,
         \ab[14][17] , \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] ,
         \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] ,
         \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] ,
         \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][21] , \ab[13][20] ,
         \ab[13][19] , \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] ,
         \ab[13][14] , \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] ,
         \ab[13][9] , \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] ,
         \ab[13][4] , \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] ,
         \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] , \ab[12][17] ,
         \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] ,
         \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] ,
         \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] ,
         \ab[12][1] , \ab[12][0] , \ab[11][21] , \ab[11][20] , \ab[11][19] ,
         \ab[11][18] , \ab[11][17] , \ab[11][16] , \ab[11][15] , \ab[11][14] ,
         \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] ,
         \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][21] ,
         \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][21] , \ab[9][20] , \ab[9][19] , \ab[9][18] ,
         \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] ,
         \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] ,
         \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] ,
         \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][21] , \ab[8][20] ,
         \ab[8][19] , \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] ,
         \ab[8][14] , \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] ,
         \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] ,
         \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][21] , \ab[6][20] , \ab[6][19] ,
         \ab[6][18] , \ab[6][17] , \ab[6][16] , \ab[6][15] , \ab[6][14] ,
         \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] ,
         \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][21] , \ab[4][20] , \ab[4][19] , \ab[4][18] ,
         \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] ,
         \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][21] , \ab[1][20] , \ab[1][19] ,
         \ab[1][18] , \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] ,
         \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] ,
         \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[24][15] ,
         \CARRYB[24][14] , \CARRYB[24][13] , \CARRYB[24][12] ,
         \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] , \CARRYB[24][8] ,
         \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] ,
         \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][20] , \CARRYB[23][19] , \CARRYB[23][18] ,
         \CARRYB[23][17] , \CARRYB[23][16] , \CARRYB[23][15] ,
         \CARRYB[23][14] , \CARRYB[23][13] , \CARRYB[23][12] ,
         \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] ,
         \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] ,
         \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] ,
         \CARRYB[22][20] , \CARRYB[22][19] , \CARRYB[22][18] ,
         \CARRYB[22][17] , \CARRYB[22][16] , \CARRYB[22][15] ,
         \CARRYB[22][14] , \CARRYB[22][13] , \CARRYB[22][12] ,
         \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] ,
         \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] ,
         \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] ,
         \CARRYB[21][20] , \CARRYB[21][19] , \CARRYB[21][18] ,
         \CARRYB[21][17] , \CARRYB[21][16] , \CARRYB[21][15] ,
         \CARRYB[21][14] , \CARRYB[21][13] , \CARRYB[21][12] ,
         \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] ,
         \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] ,
         \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] ,
         \CARRYB[20][20] , \CARRYB[20][19] , \CARRYB[20][18] ,
         \CARRYB[20][17] , \CARRYB[20][16] , \CARRYB[20][15] ,
         \CARRYB[20][14] , \CARRYB[20][13] , \CARRYB[20][12] ,
         \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] ,
         \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][20] , \CARRYB[19][19] , \CARRYB[19][18] ,
         \CARRYB[19][17] , \CARRYB[19][16] , \CARRYB[19][15] ,
         \CARRYB[19][14] , \CARRYB[19][13] , \CARRYB[19][12] ,
         \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] ,
         \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] ,
         \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] ,
         \CARRYB[18][20] , \CARRYB[18][19] , \CARRYB[18][18] ,
         \CARRYB[18][17] , \CARRYB[18][16] , \CARRYB[18][15] ,
         \CARRYB[18][14] , \CARRYB[18][13] , \CARRYB[18][12] ,
         \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] , \CARRYB[18][8] ,
         \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] , \CARRYB[18][4] ,
         \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] ,
         \CARRYB[17][20] , \CARRYB[17][19] , \CARRYB[17][18] ,
         \CARRYB[17][17] , \CARRYB[17][16] , \CARRYB[17][15] ,
         \CARRYB[17][14] , \CARRYB[17][13] , \CARRYB[17][12] ,
         \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] ,
         \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] ,
         \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] ,
         \CARRYB[16][20] , \CARRYB[16][19] , \CARRYB[16][18] ,
         \CARRYB[16][17] , \CARRYB[16][16] , \CARRYB[16][15] ,
         \CARRYB[16][14] , \CARRYB[16][13] , \CARRYB[16][12] ,
         \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] ,
         \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] ,
         \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] ,
         \CARRYB[15][20] , \CARRYB[15][19] , \CARRYB[15][18] ,
         \CARRYB[15][17] , \CARRYB[15][16] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][20] , \CARRYB[14][19] , \CARRYB[14][18] ,
         \CARRYB[14][17] , \CARRYB[14][16] , \CARRYB[14][15] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][20] , \CARRYB[13][19] , \CARRYB[13][18] ,
         \CARRYB[13][17] , \CARRYB[13][16] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][20] , \CARRYB[12][19] , \CARRYB[12][18] ,
         \CARRYB[12][17] , \CARRYB[12][16] , \CARRYB[12][15] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][20] , \CARRYB[11][19] , \CARRYB[11][18] ,
         \CARRYB[11][17] , \CARRYB[11][16] , \CARRYB[11][15] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][20] , \CARRYB[10][19] , \CARRYB[10][18] ,
         \CARRYB[10][17] , \CARRYB[10][16] , \CARRYB[10][15] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] ,
         \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] ,
         \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][20] , \CARRYB[7][19] ,
         \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] ,
         \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] ,
         \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][20] ,
         \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] ,
         \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] ,
         \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] ,
         \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][20] , \CARRYB[3][19] ,
         \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] ,
         \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][20] ,
         \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] ,
         \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] ,
         \SUMB[24][12] , \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] ,
         \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] ,
         \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] ,
         \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] ,
         \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] ,
         \SUMB[23][12] , \SUMB[23][11] , \SUMB[23][10] , \SUMB[23][9] ,
         \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] ,
         \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] ,
         \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] ,
         \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] ,
         \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] ,
         \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] ,
         \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] ,
         \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] ,
         \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] ,
         \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] ,
         \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] ,
         \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] ,
         \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] ,
         \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] ,
         \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] ,
         \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] ,
         \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][20] , \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] ,
         \SUMB[16][16] , \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] ,
         \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] ,
         \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] , \SUMB[14][17] ,
         \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] ,
         \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] ,
         \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] ,
         \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] ,
         \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] ,
         \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] ,
         \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][20] ,
         \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] ,
         \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] ,
         \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] ,
         \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][20] ,
         \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][20] ,
         \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] , \SUMB[2][16] ,
         \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] ,
         \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] ,
         \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] ,
         \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][20] , \SUMB[1][19] ,
         \SUMB[1][18] , \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] ,
         \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \PROD1[21] , \CARRYB[47][20] , \CARRYB[47][19] , \CARRYB[47][18] ,
         \CARRYB[47][17] , \CARRYB[47][16] , \CARRYB[47][15] ,
         \CARRYB[47][14] , \CARRYB[47][13] , \CARRYB[47][12] ,
         \CARRYB[47][11] , \CARRYB[47][10] , \CARRYB[47][9] , \CARRYB[47][8] ,
         \CARRYB[47][7] , \CARRYB[47][6] , \CARRYB[47][5] , \CARRYB[47][4] ,
         \CARRYB[47][3] , \CARRYB[47][2] , \CARRYB[47][1] , \CARRYB[47][0] ,
         \CARRYB[46][20] , \CARRYB[46][19] , \CARRYB[46][18] ,
         \CARRYB[46][17] , \CARRYB[46][16] , \CARRYB[46][15] ,
         \CARRYB[46][14] , \CARRYB[46][13] , \CARRYB[46][12] ,
         \CARRYB[46][11] , \CARRYB[46][10] , \CARRYB[46][9] , \CARRYB[46][8] ,
         \CARRYB[46][7] , \CARRYB[46][6] , \CARRYB[46][5] , \CARRYB[46][4] ,
         \CARRYB[46][3] , \CARRYB[46][2] , \CARRYB[46][1] , \CARRYB[46][0] ,
         \CARRYB[45][20] , \CARRYB[45][19] , \CARRYB[45][18] ,
         \CARRYB[45][17] , \CARRYB[45][16] , \CARRYB[45][15] ,
         \CARRYB[45][14] , \CARRYB[45][13] , \CARRYB[45][12] ,
         \CARRYB[45][11] , \CARRYB[45][10] , \CARRYB[45][9] , \CARRYB[45][8] ,
         \CARRYB[45][7] , \CARRYB[45][6] , \CARRYB[45][5] , \CARRYB[45][4] ,
         \CARRYB[45][3] , \CARRYB[45][2] , \CARRYB[45][1] , \CARRYB[45][0] ,
         \CARRYB[44][20] , \CARRYB[44][19] , \CARRYB[44][18] ,
         \CARRYB[44][17] , \CARRYB[44][16] , \CARRYB[44][15] ,
         \CARRYB[44][14] , \CARRYB[44][13] , \CARRYB[44][12] ,
         \CARRYB[44][11] , \CARRYB[44][10] , \CARRYB[44][9] , \CARRYB[44][8] ,
         \CARRYB[44][7] , \CARRYB[44][6] , \CARRYB[44][5] , \CARRYB[44][4] ,
         \CARRYB[44][3] , \CARRYB[44][2] , \CARRYB[44][1] , \CARRYB[44][0] ,
         \CARRYB[43][20] , \CARRYB[43][19] , \CARRYB[43][18] ,
         \CARRYB[43][17] , \CARRYB[43][16] , \CARRYB[43][15] ,
         \CARRYB[43][14] , \CARRYB[43][13] , \CARRYB[43][12] ,
         \CARRYB[43][11] , \CARRYB[43][10] , \CARRYB[43][9] , \CARRYB[43][8] ,
         \CARRYB[43][7] , \CARRYB[43][6] , \CARRYB[43][5] , \CARRYB[43][4] ,
         \CARRYB[43][3] , \CARRYB[43][2] , \CARRYB[43][1] , \CARRYB[43][0] ,
         \CARRYB[42][20] , \CARRYB[42][19] , \CARRYB[42][18] ,
         \CARRYB[42][17] , \CARRYB[42][16] , \CARRYB[42][15] ,
         \CARRYB[42][14] , \CARRYB[42][13] , \CARRYB[42][12] ,
         \CARRYB[42][11] , \CARRYB[42][10] , \CARRYB[42][9] , \CARRYB[42][8] ,
         \CARRYB[42][7] , \CARRYB[42][6] , \CARRYB[42][5] , \CARRYB[42][4] ,
         \CARRYB[42][3] , \CARRYB[42][2] , \CARRYB[42][1] , \CARRYB[42][0] ,
         \CARRYB[41][20] , \CARRYB[41][19] , \CARRYB[41][18] ,
         \CARRYB[41][17] , \CARRYB[41][16] , \CARRYB[41][15] ,
         \CARRYB[41][14] , \CARRYB[41][13] , \CARRYB[41][12] ,
         \CARRYB[41][11] , \CARRYB[41][10] , \CARRYB[41][9] , \CARRYB[41][8] ,
         \CARRYB[41][7] , \CARRYB[41][6] , \CARRYB[41][5] , \CARRYB[41][4] ,
         \CARRYB[41][3] , \CARRYB[41][2] , \CARRYB[41][1] , \CARRYB[41][0] ,
         \CARRYB[40][20] , \CARRYB[40][19] , \CARRYB[40][18] ,
         \CARRYB[40][17] , \CARRYB[40][16] , \CARRYB[40][15] ,
         \CARRYB[40][14] , \CARRYB[40][13] , \CARRYB[40][12] ,
         \CARRYB[40][11] , \CARRYB[40][10] , \CARRYB[40][9] , \CARRYB[40][8] ,
         \CARRYB[40][7] , \CARRYB[40][6] , \CARRYB[40][5] , \CARRYB[40][4] ,
         \CARRYB[40][3] , \CARRYB[40][2] , \CARRYB[40][1] , \CARRYB[40][0] ,
         \CARRYB[39][20] , \CARRYB[39][19] , \CARRYB[39][18] ,
         \CARRYB[39][17] , \CARRYB[39][16] , \CARRYB[39][15] ,
         \CARRYB[39][14] , \CARRYB[39][13] , \CARRYB[39][12] ,
         \CARRYB[39][11] , \CARRYB[39][10] , \CARRYB[39][9] , \CARRYB[39][8] ,
         \CARRYB[39][7] , \CARRYB[39][6] , \CARRYB[39][5] , \CARRYB[39][4] ,
         \CARRYB[39][3] , \CARRYB[39][2] , \CARRYB[39][1] , \CARRYB[39][0] ,
         \CARRYB[38][20] , \CARRYB[38][19] , \CARRYB[38][18] ,
         \CARRYB[38][17] , \CARRYB[38][16] , \CARRYB[38][15] ,
         \CARRYB[38][14] , \CARRYB[38][13] , \CARRYB[38][12] ,
         \CARRYB[38][11] , \CARRYB[38][10] , \CARRYB[38][9] , \CARRYB[38][8] ,
         \CARRYB[38][7] , \CARRYB[38][6] , \CARRYB[38][5] , \CARRYB[38][4] ,
         \CARRYB[38][3] , \CARRYB[38][2] , \CARRYB[38][1] , \CARRYB[38][0] ,
         \CARRYB[37][20] , \CARRYB[37][19] , \CARRYB[37][18] ,
         \CARRYB[37][17] , \CARRYB[37][16] , \CARRYB[37][15] ,
         \CARRYB[37][14] , \CARRYB[37][13] , \CARRYB[37][12] ,
         \CARRYB[37][11] , \CARRYB[37][10] , \CARRYB[37][9] , \CARRYB[37][8] ,
         \CARRYB[37][7] , \CARRYB[37][6] , \CARRYB[37][5] , \CARRYB[37][4] ,
         \CARRYB[37][3] , \CARRYB[37][2] , \CARRYB[37][1] , \CARRYB[37][0] ,
         \CARRYB[36][20] , \CARRYB[36][19] , \CARRYB[36][18] ,
         \CARRYB[36][17] , \CARRYB[36][16] , \CARRYB[36][15] ,
         \CARRYB[36][14] , \CARRYB[36][13] , \CARRYB[36][12] ,
         \CARRYB[36][11] , \CARRYB[36][10] , \CARRYB[36][9] , \CARRYB[36][8] ,
         \CARRYB[36][7] , \CARRYB[36][6] , \CARRYB[36][5] , \CARRYB[36][4] ,
         \CARRYB[36][3] , \CARRYB[36][2] , \CARRYB[36][1] , \CARRYB[36][0] ,
         \CARRYB[35][20] , \CARRYB[35][19] , \CARRYB[35][18] ,
         \CARRYB[35][17] , \CARRYB[35][16] , \CARRYB[35][15] ,
         \CARRYB[35][14] , \CARRYB[35][13] , \CARRYB[35][12] ,
         \CARRYB[35][11] , \CARRYB[35][10] , \CARRYB[35][9] , \CARRYB[35][8] ,
         \CARRYB[35][7] , \CARRYB[35][6] , \CARRYB[35][5] , \CARRYB[35][4] ,
         \CARRYB[35][3] , \CARRYB[35][2] , \CARRYB[35][1] , \CARRYB[35][0] ,
         \CARRYB[34][20] , \CARRYB[34][19] , \CARRYB[34][18] ,
         \CARRYB[34][17] , \CARRYB[34][16] , \CARRYB[34][15] ,
         \CARRYB[34][14] , \CARRYB[34][13] , \CARRYB[34][12] ,
         \CARRYB[34][11] , \CARRYB[34][10] , \CARRYB[34][9] , \CARRYB[34][8] ,
         \CARRYB[34][7] , \CARRYB[34][6] , \CARRYB[34][5] , \CARRYB[34][4] ,
         \CARRYB[34][3] , \CARRYB[34][2] , \CARRYB[34][1] , \CARRYB[34][0] ,
         \CARRYB[33][20] , \CARRYB[33][19] , \CARRYB[33][18] ,
         \CARRYB[33][17] , \CARRYB[33][16] , \CARRYB[33][15] ,
         \CARRYB[33][14] , \CARRYB[33][13] , \CARRYB[33][12] ,
         \CARRYB[33][11] , \CARRYB[33][10] , \CARRYB[33][9] , \CARRYB[33][8] ,
         \CARRYB[33][7] , \CARRYB[33][6] , \CARRYB[33][5] , \CARRYB[33][4] ,
         \CARRYB[33][3] , \CARRYB[33][2] , \CARRYB[33][1] , \CARRYB[33][0] ,
         \CARRYB[32][20] , \CARRYB[32][19] , \CARRYB[32][18] ,
         \CARRYB[32][17] , \CARRYB[32][16] , \CARRYB[32][15] ,
         \CARRYB[32][14] , \CARRYB[32][13] , \CARRYB[32][12] ,
         \CARRYB[32][11] , \CARRYB[32][10] , \CARRYB[32][9] , \CARRYB[32][8] ,
         \CARRYB[32][7] , \CARRYB[32][6] , \CARRYB[32][5] , \CARRYB[32][4] ,
         \CARRYB[32][3] , \CARRYB[32][2] , \CARRYB[32][1] , \CARRYB[32][0] ,
         \CARRYB[31][20] , \CARRYB[31][19] , \CARRYB[31][18] ,
         \CARRYB[31][17] , \CARRYB[31][16] , \CARRYB[31][15] ,
         \CARRYB[31][14] , \CARRYB[31][13] , \CARRYB[31][12] ,
         \CARRYB[31][11] , \CARRYB[31][10] , \CARRYB[31][9] , \CARRYB[31][8] ,
         \CARRYB[31][7] , \CARRYB[31][6] , \CARRYB[31][5] , \CARRYB[31][4] ,
         \CARRYB[31][3] , \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] ,
         \CARRYB[30][20] , \CARRYB[30][19] , \CARRYB[30][18] ,
         \CARRYB[30][17] , \CARRYB[30][16] , \CARRYB[30][15] ,
         \CARRYB[30][14] , \CARRYB[30][13] , \CARRYB[30][12] ,
         \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] ,
         \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] ,
         \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] ,
         \CARRYB[29][20] , \CARRYB[29][19] , \CARRYB[29][18] ,
         \CARRYB[29][17] , \CARRYB[29][16] , \CARRYB[29][15] ,
         \CARRYB[29][14] , \CARRYB[29][13] , \CARRYB[29][12] ,
         \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] , \CARRYB[29][8] ,
         \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] , \CARRYB[29][4] ,
         \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] , \CARRYB[29][0] ,
         \CARRYB[28][20] , \CARRYB[28][19] , \CARRYB[28][18] ,
         \CARRYB[28][17] , \CARRYB[28][16] , \CARRYB[28][15] ,
         \CARRYB[28][14] , \CARRYB[28][13] , \CARRYB[28][12] ,
         \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] , \CARRYB[28][8] ,
         \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] , \CARRYB[28][4] ,
         \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] ,
         \CARRYB[27][20] , \CARRYB[27][19] , \CARRYB[27][18] ,
         \CARRYB[27][17] , \CARRYB[27][16] , \CARRYB[27][15] ,
         \CARRYB[27][14] , \CARRYB[27][13] , \CARRYB[27][12] ,
         \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] , \CARRYB[27][8] ,
         \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] , \CARRYB[27][4] ,
         \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] ,
         \CARRYB[26][20] , \CARRYB[26][19] , \CARRYB[26][18] ,
         \CARRYB[26][17] , \CARRYB[26][16] , \CARRYB[26][15] ,
         \CARRYB[26][14] , \CARRYB[26][13] , \CARRYB[26][12] ,
         \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] , \CARRYB[26][8] ,
         \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] , \CARRYB[26][4] ,
         \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] , \CARRYB[26][0] ,
         \CARRYB[25][20] , \CARRYB[25][19] , \CARRYB[25][18] ,
         \CARRYB[25][17] , \CARRYB[25][16] , \CARRYB[25][15] ,
         \CARRYB[25][14] , \CARRYB[25][13] , \CARRYB[25][12] ,
         \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][9] , \CARRYB[25][8] ,
         \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] ,
         \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] ,
         \CARRYB[24][20] , \CARRYB[24][19] , \CARRYB[24][18] ,
         \CARRYB[24][17] , \CARRYB[24][16] , \SUMB[47][20] , \SUMB[47][19] ,
         \SUMB[47][18] , \SUMB[47][17] , \SUMB[47][16] , \SUMB[47][15] ,
         \SUMB[47][14] , \SUMB[47][13] , \SUMB[47][12] , \SUMB[47][11] ,
         \SUMB[47][10] , \SUMB[47][9] , \SUMB[47][8] , \SUMB[47][7] ,
         \SUMB[47][6] , \SUMB[47][5] , \SUMB[47][4] , \SUMB[47][3] ,
         \SUMB[47][2] , \SUMB[47][1] , \SUMB[47][0] , \SUMB[46][20] ,
         \SUMB[46][19] , \SUMB[46][18] , \SUMB[46][17] , \SUMB[46][16] ,
         \SUMB[46][15] , \SUMB[46][14] , \SUMB[46][13] , \SUMB[46][12] ,
         \SUMB[46][11] , \SUMB[46][10] , \SUMB[46][9] , \SUMB[46][8] ,
         \SUMB[46][7] , \SUMB[46][6] , \SUMB[46][5] , \SUMB[46][4] ,
         \SUMB[46][3] , \SUMB[46][2] , \SUMB[46][1] , \SUMB[45][20] ,
         \SUMB[45][19] , \SUMB[45][18] , \SUMB[45][17] , \SUMB[45][16] ,
         \SUMB[45][15] , \SUMB[45][14] , \SUMB[45][13] , \SUMB[45][12] ,
         \SUMB[45][11] , \SUMB[45][10] , \SUMB[45][9] , \SUMB[45][8] ,
         \SUMB[45][7] , \SUMB[45][6] , \SUMB[45][5] , \SUMB[45][4] ,
         \SUMB[45][3] , \SUMB[45][2] , \SUMB[45][1] , \SUMB[44][20] ,
         \SUMB[44][19] , \SUMB[44][18] , \SUMB[44][17] , \SUMB[44][16] ,
         \SUMB[44][15] , \SUMB[44][14] , \SUMB[44][13] , \SUMB[44][12] ,
         \SUMB[44][11] , \SUMB[44][10] , \SUMB[44][9] , \SUMB[44][8] ,
         \SUMB[44][7] , \SUMB[44][6] , \SUMB[44][5] , \SUMB[44][4] ,
         \SUMB[44][3] , \SUMB[44][2] , \SUMB[44][1] , \SUMB[43][20] ,
         \SUMB[43][19] , \SUMB[43][18] , \SUMB[43][17] , \SUMB[43][16] ,
         \SUMB[43][15] , \SUMB[43][14] , \SUMB[43][13] , \SUMB[43][12] ,
         \SUMB[43][11] , \SUMB[43][10] , \SUMB[43][9] , \SUMB[43][8] ,
         \SUMB[43][7] , \SUMB[43][6] , \SUMB[43][5] , \SUMB[43][4] ,
         \SUMB[43][3] , \SUMB[43][2] , \SUMB[43][1] , \SUMB[42][20] ,
         \SUMB[42][19] , \SUMB[42][18] , \SUMB[42][17] , \SUMB[42][16] ,
         \SUMB[42][15] , \SUMB[42][14] , \SUMB[42][13] , \SUMB[42][12] ,
         \SUMB[42][11] , \SUMB[42][10] , \SUMB[42][9] , \SUMB[42][8] ,
         \SUMB[42][7] , \SUMB[42][6] , \SUMB[42][5] , \SUMB[42][4] ,
         \SUMB[42][3] , \SUMB[42][2] , \SUMB[42][1] , \SUMB[41][20] ,
         \SUMB[41][19] , \SUMB[41][18] , \SUMB[41][17] , \SUMB[41][16] ,
         \SUMB[41][15] , \SUMB[41][14] , \SUMB[41][13] , \SUMB[41][12] ,
         \SUMB[41][11] , \SUMB[41][10] , \SUMB[41][9] , \SUMB[41][8] ,
         \SUMB[41][7] , \SUMB[41][6] , \SUMB[41][5] , \SUMB[41][4] ,
         \SUMB[41][3] , \SUMB[41][2] , \SUMB[41][1] , \SUMB[40][20] ,
         \SUMB[40][19] , \SUMB[40][18] , \SUMB[40][17] , \SUMB[40][16] ,
         \SUMB[40][15] , \SUMB[40][14] , \SUMB[40][13] , \SUMB[40][12] ,
         \SUMB[40][11] , \SUMB[40][10] , \SUMB[40][9] , \SUMB[40][8] ,
         \SUMB[40][7] , \SUMB[40][6] , \SUMB[40][5] , \SUMB[40][4] ,
         \SUMB[40][3] , \SUMB[40][2] , \SUMB[40][1] , \SUMB[39][20] ,
         \SUMB[39][19] , \SUMB[39][18] , \SUMB[39][17] , \SUMB[39][16] ,
         \SUMB[39][15] , \SUMB[39][14] , \SUMB[39][13] , \SUMB[39][12] ,
         \SUMB[39][11] , \SUMB[39][10] , \SUMB[39][9] , \SUMB[39][8] ,
         \SUMB[39][7] , \SUMB[39][6] , \SUMB[39][5] , \SUMB[39][4] ,
         \SUMB[39][3] , \SUMB[39][2] , \SUMB[39][1] , \SUMB[38][20] ,
         \SUMB[38][19] , \SUMB[38][18] , \SUMB[38][17] , \SUMB[38][16] ,
         \SUMB[38][15] , \SUMB[38][14] , \SUMB[38][13] , \SUMB[38][12] ,
         \SUMB[38][11] , \SUMB[38][10] , \SUMB[38][9] , \SUMB[38][8] ,
         \SUMB[38][7] , \SUMB[38][6] , \SUMB[38][5] , \SUMB[38][4] ,
         \SUMB[38][3] , \SUMB[38][2] , \SUMB[38][1] , \SUMB[37][20] ,
         \SUMB[37][19] , \SUMB[37][18] , \SUMB[37][17] , \SUMB[37][16] ,
         \SUMB[37][15] , \SUMB[37][14] , \SUMB[37][13] , \SUMB[37][12] ,
         \SUMB[37][11] , \SUMB[37][10] , \SUMB[37][9] , \SUMB[37][8] ,
         \SUMB[37][7] , \SUMB[37][6] , \SUMB[37][5] , \SUMB[37][4] ,
         \SUMB[37][3] , \SUMB[37][2] , \SUMB[37][1] , \SUMB[36][20] ,
         \SUMB[36][19] , \SUMB[36][18] , \SUMB[36][17] , \SUMB[36][16] ,
         \SUMB[36][15] , \SUMB[36][14] , \SUMB[36][13] , \SUMB[36][12] ,
         \SUMB[36][11] , \SUMB[36][10] , \SUMB[36][9] , \SUMB[36][8] ,
         \SUMB[36][7] , \SUMB[36][6] , \SUMB[36][5] , \SUMB[36][4] ,
         \SUMB[36][3] , \SUMB[36][2] , \SUMB[36][1] , \SUMB[35][20] ,
         \SUMB[35][19] , \SUMB[35][18] , \SUMB[35][17] , \SUMB[35][16] ,
         \SUMB[35][15] , \SUMB[35][14] , \SUMB[35][13] , \SUMB[35][12] ,
         \SUMB[35][11] , \SUMB[35][10] , \SUMB[35][9] , \SUMB[35][8] ,
         \SUMB[35][7] , \SUMB[35][6] , \SUMB[35][5] , \SUMB[35][4] ,
         \SUMB[35][3] , \SUMB[35][2] , \SUMB[35][1] , \SUMB[34][20] ,
         \SUMB[34][19] , \SUMB[34][18] , \SUMB[34][17] , \SUMB[34][16] ,
         \SUMB[34][15] , \SUMB[34][14] , \SUMB[34][13] , \SUMB[34][12] ,
         \SUMB[34][11] , \SUMB[34][10] , \SUMB[34][9] , \SUMB[34][8] ,
         \SUMB[34][7] , \SUMB[34][6] , \SUMB[34][5] , \SUMB[34][4] ,
         \SUMB[34][3] , \SUMB[34][2] , \SUMB[34][1] , \SUMB[33][20] ,
         \SUMB[33][19] , \SUMB[33][18] , \SUMB[33][17] , \SUMB[33][16] ,
         \SUMB[33][15] , \SUMB[33][14] , \SUMB[33][13] , \SUMB[33][12] ,
         \SUMB[33][11] , \SUMB[33][10] , \SUMB[33][9] , \SUMB[33][8] ,
         \SUMB[33][7] , \SUMB[33][6] , \SUMB[33][5] , \SUMB[33][4] ,
         \SUMB[33][3] , \SUMB[33][2] , \SUMB[33][1] , \SUMB[32][20] ,
         \SUMB[32][19] , \SUMB[32][18] , \SUMB[32][17] , \SUMB[32][16] ,
         \SUMB[32][15] , \SUMB[32][14] , \SUMB[32][13] , \SUMB[32][12] ,
         \SUMB[32][11] , \SUMB[32][10] , \SUMB[32][9] , \SUMB[32][8] ,
         \SUMB[32][7] , \SUMB[32][6] , \SUMB[32][5] , \SUMB[32][4] ,
         \SUMB[32][3] , \SUMB[32][2] , \SUMB[32][1] , \SUMB[31][20] ,
         \SUMB[31][19] , \SUMB[31][18] , \SUMB[31][17] , \SUMB[31][16] ,
         \SUMB[31][15] , \SUMB[31][14] , \SUMB[31][13] , \SUMB[31][12] ,
         \SUMB[31][11] , \SUMB[31][10] , \SUMB[31][9] , \SUMB[31][8] ,
         \SUMB[31][7] , \SUMB[31][6] , \SUMB[31][5] , \SUMB[31][4] ,
         \SUMB[31][3] , \SUMB[31][2] , \SUMB[31][1] , \SUMB[30][20] ,
         \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] , \SUMB[30][16] ,
         \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] , \SUMB[30][12] ,
         \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][20] ,
         \SUMB[29][19] , \SUMB[29][18] , \SUMB[29][17] , \SUMB[29][16] ,
         \SUMB[29][15] , \SUMB[29][14] , \SUMB[29][13] , \SUMB[29][12] ,
         \SUMB[29][11] , \SUMB[29][10] , \SUMB[29][9] , \SUMB[29][8] ,
         \SUMB[29][7] , \SUMB[29][6] , \SUMB[29][5] , \SUMB[29][4] ,
         \SUMB[29][3] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][20] ,
         \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] ,
         \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] ,
         \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] ,
         \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] ,
         \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][20] ,
         \SUMB[27][19] , \SUMB[27][18] , \SUMB[27][17] , \SUMB[27][16] ,
         \SUMB[27][15] , \SUMB[27][14] , \SUMB[27][13] , \SUMB[27][12] ,
         \SUMB[27][11] , \SUMB[27][10] , \SUMB[27][9] , \SUMB[27][8] ,
         \SUMB[27][7] , \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] ,
         \SUMB[27][3] , \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][20] ,
         \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] , \SUMB[26][16] ,
         \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] , \SUMB[26][12] ,
         \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] , \SUMB[26][8] ,
         \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][20] ,
         \SUMB[25][19] , \SUMB[25][18] , \SUMB[25][17] , \SUMB[25][16] ,
         \SUMB[25][15] , \SUMB[25][14] , \SUMB[25][13] , \SUMB[25][12] ,
         \SUMB[25][11] , \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] ,
         \SUMB[25][7] , \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] ,
         \SUMB[25][3] , \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][20] ,
         \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] , \SUMB[24][16] ,
         \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] ,
         \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] ,
         \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] ,
         \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] ,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[18] , \A1[17] , \A1[16] ,
         \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] ,
         \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] ,
         \A1[1] , \A1[0] , \A2[67] , \A2[66] , \A2[65] , \A2[64] , \A2[63] ,
         \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] ,
         \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] ,
         \A2[48] , \A2[47] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37;

  Poly_Logarithm_DW01_add_2 FS_1 ( .A({1'b0, \A1[66] , \A1[65] , \A1[64] , 
        \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , 
        \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , 
        \A1[49] , \A1[48] , \A1[47] , \A1[46] , \SUMB[47][0] , \A1[44] , 
        \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , 
        \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , 
        \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , 
        \A1[22] , \A1[21] , \A1[20] , \PROD1[21] , \A1[18] , \A1[17] , 
        \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({\A2[67] , \A2[66] , \A2[65] , \A2[64] , 
        \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , 
        \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , 
        \A2[49] , \A2[48] , \A2[47] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, PRODUCT[67:38], SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S4_0 ( .A(\ab[47][0] ), .B(\CARRYB[46][0] ), .CI(\SUMB[46][1] ), .CO(
        \CARRYB[47][0] ), .S(\SUMB[47][0] ) );
  FA1A S1_46_0 ( .A(\ab[46][0] ), .B(\CARRYB[45][0] ), .CI(\SUMB[45][1] ), 
        .CO(\CARRYB[46][0] ), .S(\A1[44] ) );
  FA1A S1_45_0 ( .A(\ab[45][0] ), .B(\CARRYB[44][0] ), .CI(\SUMB[44][1] ), 
        .CO(\CARRYB[45][0] ), .S(\A1[43] ) );
  FA1A S1_44_0 ( .A(\ab[44][0] ), .B(\CARRYB[43][0] ), .CI(\SUMB[43][1] ), 
        .CO(\CARRYB[44][0] ), .S(\A1[42] ) );
  FA1A S1_43_0 ( .A(\ab[43][0] ), .B(\CARRYB[42][0] ), .CI(\SUMB[42][1] ), 
        .CO(\CARRYB[43][0] ), .S(\A1[41] ) );
  FA1A S1_42_0 ( .A(\ab[42][0] ), .B(\CARRYB[41][0] ), .CI(\SUMB[41][1] ), 
        .CO(\CARRYB[42][0] ), .S(\A1[40] ) );
  FA1A S1_41_0 ( .A(\ab[41][0] ), .B(\CARRYB[40][0] ), .CI(\SUMB[40][1] ), 
        .CO(\CARRYB[41][0] ), .S(\A1[39] ) );
  FA1A S1_40_0 ( .A(\ab[40][0] ), .B(\CARRYB[39][0] ), .CI(\SUMB[39][1] ), 
        .CO(\CARRYB[40][0] ), .S(\A1[38] ) );
  FA1A S1_39_0 ( .A(\ab[39][0] ), .B(\CARRYB[38][0] ), .CI(\SUMB[38][1] ), 
        .CO(\CARRYB[39][0] ), .S(\A1[37] ) );
  FA1A S1_36_0 ( .A(\ab[36][0] ), .B(\CARRYB[35][0] ), .CI(\SUMB[35][1] ), 
        .CO(\CARRYB[36][0] ), .S(\A1[34] ) );
  FA1A S1_37_0 ( .A(\ab[37][0] ), .B(\CARRYB[36][0] ), .CI(\SUMB[36][1] ), 
        .CO(\CARRYB[37][0] ), .S(\A1[35] ) );
  FA1A S1_38_0 ( .A(\ab[38][0] ), .B(\CARRYB[37][0] ), .CI(\SUMB[37][1] ), 
        .CO(\CARRYB[38][0] ), .S(\A1[36] ) );
  FA1A S5_20 ( .A(\ab[47][20] ), .B(\CARRYB[46][20] ), .CI(\ab[46][21] ), .CO(
        \CARRYB[47][20] ), .S(\SUMB[47][20] ) );
  FA1A S4_19 ( .A(\ab[47][19] ), .B(\CARRYB[46][19] ), .CI(\SUMB[46][20] ), 
        .CO(\CARRYB[47][19] ), .S(\SUMB[47][19] ) );
  FA1A S3_46_20 ( .A(\ab[46][20] ), .B(\CARRYB[45][20] ), .CI(\ab[45][21] ), 
        .CO(\CARRYB[46][20] ), .S(\SUMB[46][20] ) );
  FA1A S2_36_1 ( .A(\ab[36][1] ), .B(\CARRYB[35][1] ), .CI(\SUMB[35][2] ), 
        .CO(\CARRYB[36][1] ), .S(\SUMB[36][1] ) );
  FA1A S4_18 ( .A(\ab[47][18] ), .B(\CARRYB[46][18] ), .CI(\SUMB[46][19] ), 
        .CO(\CARRYB[47][18] ), .S(\SUMB[47][18] ) );
  FA1A S1_33_0 ( .A(\ab[33][0] ), .B(\CARRYB[32][0] ), .CI(\SUMB[32][1] ), 
        .CO(\CARRYB[33][0] ), .S(\A1[31] ) );
  FA1A S1_34_0 ( .A(\ab[34][0] ), .B(\CARRYB[33][0] ), .CI(\SUMB[33][1] ), 
        .CO(\CARRYB[34][0] ), .S(\A1[32] ) );
  FA1A S1_35_0 ( .A(\ab[35][0] ), .B(\CARRYB[34][0] ), .CI(\SUMB[34][1] ), 
        .CO(\CARRYB[35][0] ), .S(\A1[33] ) );
  FA1A S2_35_1 ( .A(\ab[35][1] ), .B(\CARRYB[34][1] ), .CI(\SUMB[34][2] ), 
        .CO(\CARRYB[35][1] ), .S(\SUMB[35][1] ) );
  FA1A S2_46_19 ( .A(\ab[46][19] ), .B(\CARRYB[45][19] ), .CI(\SUMB[45][20] ), 
        .CO(\CARRYB[46][19] ), .S(\SUMB[46][19] ) );
  FA1A S2_34_1 ( .A(\ab[34][1] ), .B(\CARRYB[33][1] ), .CI(\SUMB[33][2] ), 
        .CO(\CARRYB[34][1] ), .S(\SUMB[34][1] ) );
  FA1A S3_45_20 ( .A(\ab[45][20] ), .B(\CARRYB[44][20] ), .CI(\ab[44][21] ), 
        .CO(\CARRYB[45][20] ), .S(\SUMB[45][20] ) );
  FA1A S4_16 ( .A(\ab[47][16] ), .B(\CARRYB[46][16] ), .CI(\SUMB[46][17] ), 
        .CO(\CARRYB[47][16] ), .S(\SUMB[47][16] ) );
  FA1A S4_17 ( .A(\ab[47][17] ), .B(\CARRYB[46][17] ), .CI(\SUMB[46][18] ), 
        .CO(\CARRYB[47][17] ), .S(\SUMB[47][17] ) );
  FA1A S4_15 ( .A(\ab[47][15] ), .B(\CARRYB[46][15] ), .CI(\SUMB[46][16] ), 
        .CO(\CARRYB[47][15] ), .S(\SUMB[47][15] ) );
  FA1A S4_2 ( .A(\ab[47][2] ), .B(\CARRYB[46][2] ), .CI(\SUMB[46][3] ), .CO(
        \CARRYB[47][2] ), .S(\SUMB[47][2] ) );
  FA1A S2_33_1 ( .A(\ab[33][1] ), .B(\CARRYB[32][1] ), .CI(\SUMB[32][2] ), 
        .CO(\CARRYB[33][1] ), .S(\SUMB[33][1] ) );
  FA1A S2_46_16 ( .A(\ab[46][16] ), .B(\CARRYB[45][16] ), .CI(\SUMB[45][17] ), 
        .CO(\CARRYB[46][16] ), .S(\SUMB[46][16] ) );
  FA1A S2_46_17 ( .A(\ab[46][17] ), .B(\CARRYB[45][17] ), .CI(\SUMB[45][18] ), 
        .CO(\CARRYB[46][17] ), .S(\SUMB[46][17] ) );
  FA1A S2_46_18 ( .A(\ab[46][18] ), .B(\CARRYB[45][18] ), .CI(\SUMB[45][19] ), 
        .CO(\CARRYB[46][18] ), .S(\SUMB[46][18] ) );
  FA1A S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(\A1[28] ) );
  FA1A S1_31_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), 
        .CO(\CARRYB[31][0] ), .S(\A1[29] ) );
  FA1A S1_32_0 ( .A(\ab[32][0] ), .B(\CARRYB[31][0] ), .CI(\SUMB[31][1] ), 
        .CO(\CARRYB[32][0] ), .S(\A1[30] ) );
  FA1A S2_32_1 ( .A(\ab[32][1] ), .B(\CARRYB[31][1] ), .CI(\SUMB[31][2] ), 
        .CO(\CARRYB[32][1] ), .S(\SUMB[32][1] ) );
  FA1A S2_45_17 ( .A(\ab[45][17] ), .B(\CARRYB[44][17] ), .CI(\SUMB[44][18] ), 
        .CO(\CARRYB[45][17] ), .S(\SUMB[45][17] ) );
  FA1A S2_45_18 ( .A(\ab[45][18] ), .B(\CARRYB[44][18] ), .CI(\SUMB[44][19] ), 
        .CO(\CARRYB[45][18] ), .S(\SUMB[45][18] ) );
  FA1A S2_45_19 ( .A(\ab[45][19] ), .B(\CARRYB[44][19] ), .CI(\SUMB[44][20] ), 
        .CO(\CARRYB[45][19] ), .S(\SUMB[45][19] ) );
  FA1A S2_31_1 ( .A(\ab[31][1] ), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), 
        .CO(\CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FA1A S2_44_18 ( .A(\ab[44][18] ), .B(\CARRYB[43][18] ), .CI(\SUMB[43][19] ), 
        .CO(\CARRYB[44][18] ), .S(\SUMB[44][18] ) );
  FA1A S2_44_19 ( .A(\ab[44][19] ), .B(\CARRYB[43][19] ), .CI(\SUMB[43][20] ), 
        .CO(\CARRYB[44][19] ), .S(\SUMB[44][19] ) );
  FA1A S3_44_20 ( .A(\ab[44][20] ), .B(\CARRYB[43][20] ), .CI(\ab[43][21] ), 
        .CO(\CARRYB[44][20] ), .S(\SUMB[44][20] ) );
  FA1A S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA1A S4_14 ( .A(\ab[47][14] ), .B(\CARRYB[46][14] ), .CI(\SUMB[46][15] ), 
        .CO(\CARRYB[47][14] ), .S(\SUMB[47][14] ) );
  FA1A S2_43_19 ( .A(\ab[43][19] ), .B(\CARRYB[42][19] ), .CI(\SUMB[42][20] ), 
        .CO(\CARRYB[43][19] ), .S(\SUMB[43][19] ) );
  FA1A S3_43_20 ( .A(\ab[43][20] ), .B(\CARRYB[42][20] ), .CI(\ab[42][21] ), 
        .CO(\CARRYB[43][20] ), .S(\SUMB[43][20] ) );
  FA1A S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA1A S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA1A S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FA1A S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1A S2_46_15 ( .A(\ab[46][15] ), .B(\CARRYB[45][15] ), .CI(\SUMB[45][16] ), 
        .CO(\CARRYB[46][15] ), .S(\SUMB[46][15] ) );
  FA1A S3_42_20 ( .A(\ab[42][20] ), .B(\CARRYB[41][20] ), .CI(\ab[41][21] ), 
        .CO(\CARRYB[42][20] ), .S(\SUMB[42][20] ) );
  FA1A S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1A S2_45_16 ( .A(\ab[45][16] ), .B(\CARRYB[44][16] ), .CI(\SUMB[44][17] ), 
        .CO(\CARRYB[45][16] ), .S(\SUMB[45][16] ) );
  FA1A S4_12 ( .A(\ab[47][12] ), .B(\CARRYB[46][12] ), .CI(\SUMB[46][13] ), 
        .CO(\CARRYB[47][12] ), .S(\SUMB[47][12] ) );
  FA1A S4_13 ( .A(\ab[47][13] ), .B(\CARRYB[46][13] ), .CI(\SUMB[46][14] ), 
        .CO(\CARRYB[47][13] ), .S(\SUMB[47][13] ) );
  FA1A S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1A S2_44_17 ( .A(\ab[44][17] ), .B(\CARRYB[43][17] ), .CI(\SUMB[43][18] ), 
        .CO(\CARRYB[44][17] ), .S(\SUMB[44][17] ) );
  FA1A S2_46_13 ( .A(\ab[46][13] ), .B(\CARRYB[45][13] ), .CI(\SUMB[45][14] ), 
        .CO(\CARRYB[46][13] ), .S(\SUMB[46][13] ) );
  FA1A S2_46_14 ( .A(\ab[46][14] ), .B(\CARRYB[45][14] ), .CI(\SUMB[45][15] ), 
        .CO(\CARRYB[46][14] ), .S(\SUMB[46][14] ) );
  FA1A S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA1A S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA1A S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA1A S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S2_43_18 ( .A(\ab[43][18] ), .B(\CARRYB[42][18] ), .CI(\SUMB[42][19] ), 
        .CO(\CARRYB[43][18] ), .S(\SUMB[43][18] ) );
  FA1A S2_45_14 ( .A(\ab[45][14] ), .B(\CARRYB[44][14] ), .CI(\SUMB[44][15] ), 
        .CO(\CARRYB[45][14] ), .S(\SUMB[45][14] ) );
  FA1A S2_45_15 ( .A(\ab[45][15] ), .B(\CARRYB[44][15] ), .CI(\SUMB[44][16] ), 
        .CO(\CARRYB[45][15] ), .S(\SUMB[45][15] ) );
  FA1A S4_8 ( .A(\ab[47][8] ), .B(\CARRYB[46][8] ), .CI(\SUMB[46][9] ), .CO(
        \CARRYB[47][8] ), .S(\SUMB[47][8] ) );
  FA1A S4_9 ( .A(\ab[47][9] ), .B(\CARRYB[46][9] ), .CI(\SUMB[46][10] ), .CO(
        \CARRYB[47][9] ), .S(\SUMB[47][9] ) );
  FA1A S4_10 ( .A(\ab[47][10] ), .B(\CARRYB[46][10] ), .CI(\SUMB[46][11] ), 
        .CO(\CARRYB[47][10] ), .S(\SUMB[47][10] ) );
  FA1A S4_6 ( .A(\ab[47][6] ), .B(\CARRYB[46][6] ), .CI(\SUMB[46][7] ), .CO(
        \CARRYB[47][6] ), .S(\SUMB[47][6] ) );
  FA1A S4_7 ( .A(\ab[47][7] ), .B(\CARRYB[46][7] ), .CI(\SUMB[46][8] ), .CO(
        \CARRYB[47][7] ), .S(\SUMB[47][7] ) );
  FA1A S4_5 ( .A(\ab[47][5] ), .B(\CARRYB[46][5] ), .CI(\SUMB[46][6] ), .CO(
        \CARRYB[47][5] ), .S(\SUMB[47][5] ) );
  FA1A S4_4 ( .A(\ab[47][4] ), .B(\CARRYB[46][4] ), .CI(\SUMB[46][5] ), .CO(
        \CARRYB[47][4] ), .S(\SUMB[47][4] ) );
  FA1A S4_1 ( .A(\ab[47][1] ), .B(\CARRYB[46][1] ), .CI(\SUMB[46][2] ), .CO(
        \CARRYB[47][1] ), .S(\SUMB[47][1] ) );
  FA1A S4_3 ( .A(\ab[47][3] ), .B(\CARRYB[46][3] ), .CI(\SUMB[46][4] ), .CO(
        \CARRYB[47][3] ), .S(\SUMB[47][3] ) );
  FA1A S4_11 ( .A(\ab[47][11] ), .B(\CARRYB[46][11] ), .CI(\SUMB[46][12] ), 
        .CO(\CARRYB[47][11] ), .S(\SUMB[47][11] ) );
  FA1A S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA1A S2_42_19 ( .A(\ab[42][19] ), .B(\CARRYB[41][19] ), .CI(\SUMB[41][20] ), 
        .CO(\CARRYB[42][19] ), .S(\SUMB[42][19] ) );
  FA1A S2_44_15 ( .A(\ab[44][15] ), .B(\CARRYB[43][15] ), .CI(\SUMB[43][16] ), 
        .CO(\CARRYB[44][15] ), .S(\SUMB[44][15] ) );
  FA1A S2_44_16 ( .A(\ab[44][16] ), .B(\CARRYB[43][16] ), .CI(\SUMB[43][17] ), 
        .CO(\CARRYB[44][16] ), .S(\SUMB[44][16] ) );
  FA1A S2_46_8 ( .A(\ab[46][8] ), .B(\CARRYB[45][8] ), .CI(\SUMB[45][9] ), 
        .CO(\CARRYB[46][8] ), .S(\SUMB[46][8] ) );
  FA1A S2_46_9 ( .A(\ab[46][9] ), .B(\CARRYB[45][9] ), .CI(\SUMB[45][10] ), 
        .CO(\CARRYB[46][9] ), .S(\SUMB[46][9] ) );
  FA1A S2_46_10 ( .A(\ab[46][10] ), .B(\CARRYB[45][10] ), .CI(\SUMB[45][11] ), 
        .CO(\CARRYB[46][10] ), .S(\SUMB[46][10] ) );
  FA1A S2_46_11 ( .A(\ab[46][11] ), .B(\CARRYB[45][11] ), .CI(\SUMB[45][12] ), 
        .CO(\CARRYB[46][11] ), .S(\SUMB[46][11] ) );
  FA1A S2_46_6 ( .A(\ab[46][6] ), .B(\CARRYB[45][6] ), .CI(\SUMB[45][7] ), 
        .CO(\CARRYB[46][6] ), .S(\SUMB[46][6] ) );
  FA1A S2_46_7 ( .A(\ab[46][7] ), .B(\CARRYB[45][7] ), .CI(\SUMB[45][8] ), 
        .CO(\CARRYB[46][7] ), .S(\SUMB[46][7] ) );
  FA1A S2_46_5 ( .A(\ab[46][5] ), .B(\CARRYB[45][5] ), .CI(\SUMB[45][6] ), 
        .CO(\CARRYB[46][5] ), .S(\SUMB[46][5] ) );
  FA1A S2_46_4 ( .A(\ab[46][4] ), .B(\CARRYB[45][4] ), .CI(\SUMB[45][5] ), 
        .CO(\CARRYB[46][4] ), .S(\SUMB[46][4] ) );
  FA1A S2_46_1 ( .A(\ab[46][1] ), .B(\CARRYB[45][1] ), .CI(\SUMB[45][2] ), 
        .CO(\CARRYB[46][1] ), .S(\SUMB[46][1] ) );
  FA1A S2_46_2 ( .A(\ab[46][2] ), .B(\CARRYB[45][2] ), .CI(\SUMB[45][3] ), 
        .CO(\CARRYB[46][2] ), .S(\SUMB[46][2] ) );
  FA1A S2_46_3 ( .A(\ab[46][3] ), .B(\CARRYB[45][3] ), .CI(\SUMB[45][4] ), 
        .CO(\CARRYB[46][3] ), .S(\SUMB[46][3] ) );
  FA1A S2_46_12 ( .A(\ab[46][12] ), .B(\CARRYB[45][12] ), .CI(\SUMB[45][13] ), 
        .CO(\CARRYB[46][12] ), .S(\SUMB[46][12] ) );
  FA1A S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA1A S3_41_20 ( .A(\ab[41][20] ), .B(\CARRYB[40][20] ), .CI(\ab[40][21] ), 
        .CO(\CARRYB[41][20] ), .S(\SUMB[41][20] ) );
  FA1A S2_43_16 ( .A(\ab[43][16] ), .B(\CARRYB[42][16] ), .CI(\SUMB[42][17] ), 
        .CO(\CARRYB[43][16] ), .S(\SUMB[43][16] ) );
  FA1A S2_43_17 ( .A(\ab[43][17] ), .B(\CARRYB[42][17] ), .CI(\SUMB[42][18] ), 
        .CO(\CARRYB[43][17] ), .S(\SUMB[43][17] ) );
  FA1A S2_45_8 ( .A(\ab[45][8] ), .B(\CARRYB[44][8] ), .CI(\SUMB[44][9] ), 
        .CO(\CARRYB[45][8] ), .S(\SUMB[45][8] ) );
  FA1A S2_45_9 ( .A(\ab[45][9] ), .B(\CARRYB[44][9] ), .CI(\SUMB[44][10] ), 
        .CO(\CARRYB[45][9] ), .S(\SUMB[45][9] ) );
  FA1A S2_45_10 ( .A(\ab[45][10] ), .B(\CARRYB[44][10] ), .CI(\SUMB[44][11] ), 
        .CO(\CARRYB[45][10] ), .S(\SUMB[45][10] ) );
  FA1A S2_45_11 ( .A(\ab[45][11] ), .B(\CARRYB[44][11] ), .CI(\SUMB[44][12] ), 
        .CO(\CARRYB[45][11] ), .S(\SUMB[45][11] ) );
  FA1A S2_45_12 ( .A(\ab[45][12] ), .B(\CARRYB[44][12] ), .CI(\SUMB[44][13] ), 
        .CO(\CARRYB[45][12] ), .S(\SUMB[45][12] ) );
  FA1A S2_45_6 ( .A(\ab[45][6] ), .B(\CARRYB[44][6] ), .CI(\SUMB[44][7] ), 
        .CO(\CARRYB[45][6] ), .S(\SUMB[45][6] ) );
  FA1A S2_45_7 ( .A(\ab[45][7] ), .B(\CARRYB[44][7] ), .CI(\SUMB[44][8] ), 
        .CO(\CARRYB[45][7] ), .S(\SUMB[45][7] ) );
  FA1A S2_45_5 ( .A(\ab[45][5] ), .B(\CARRYB[44][5] ), .CI(\SUMB[44][6] ), 
        .CO(\CARRYB[45][5] ), .S(\SUMB[45][5] ) );
  FA1A S2_45_4 ( .A(\ab[45][4] ), .B(\CARRYB[44][4] ), .CI(\SUMB[44][5] ), 
        .CO(\CARRYB[45][4] ), .S(\SUMB[45][4] ) );
  FA1A S2_45_1 ( .A(\ab[45][1] ), .B(\CARRYB[44][1] ), .CI(\SUMB[44][2] ), 
        .CO(\CARRYB[45][1] ), .S(\SUMB[45][1] ) );
  FA1A S2_45_2 ( .A(\ab[45][2] ), .B(\CARRYB[44][2] ), .CI(\SUMB[44][3] ), 
        .CO(\CARRYB[45][2] ), .S(\SUMB[45][2] ) );
  FA1A S2_45_3 ( .A(\ab[45][3] ), .B(\CARRYB[44][3] ), .CI(\SUMB[44][4] ), 
        .CO(\CARRYB[45][3] ), .S(\SUMB[45][3] ) );
  FA1A S2_45_13 ( .A(\ab[45][13] ), .B(\CARRYB[44][13] ), .CI(\SUMB[44][14] ), 
        .CO(\CARRYB[45][13] ), .S(\SUMB[45][13] ) );
  FA1A S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\PROD1[21] ) );
  FA1A S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA1A S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA1A S2_42_17 ( .A(\ab[42][17] ), .B(\CARRYB[41][17] ), .CI(\SUMB[41][18] ), 
        .CO(\CARRYB[42][17] ), .S(\SUMB[42][17] ) );
  FA1A S2_42_18 ( .A(\ab[42][18] ), .B(\CARRYB[41][18] ), .CI(\SUMB[41][19] ), 
        .CO(\CARRYB[42][18] ), .S(\SUMB[42][18] ) );
  FA1A S2_44_8 ( .A(\ab[44][8] ), .B(\CARRYB[43][8] ), .CI(\SUMB[43][9] ), 
        .CO(\CARRYB[44][8] ), .S(\SUMB[44][8] ) );
  FA1A S2_44_9 ( .A(\ab[44][9] ), .B(\CARRYB[43][9] ), .CI(\SUMB[43][10] ), 
        .CO(\CARRYB[44][9] ), .S(\SUMB[44][9] ) );
  FA1A S2_44_10 ( .A(\ab[44][10] ), .B(\CARRYB[43][10] ), .CI(\SUMB[43][11] ), 
        .CO(\CARRYB[44][10] ), .S(\SUMB[44][10] ) );
  FA1A S2_44_11 ( .A(\ab[44][11] ), .B(\CARRYB[43][11] ), .CI(\SUMB[43][12] ), 
        .CO(\CARRYB[44][11] ), .S(\SUMB[44][11] ) );
  FA1A S2_44_12 ( .A(\ab[44][12] ), .B(\CARRYB[43][12] ), .CI(\SUMB[43][13] ), 
        .CO(\CARRYB[44][12] ), .S(\SUMB[44][12] ) );
  FA1A S2_44_13 ( .A(\ab[44][13] ), .B(\CARRYB[43][13] ), .CI(\SUMB[43][14] ), 
        .CO(\CARRYB[44][13] ), .S(\SUMB[44][13] ) );
  FA1A S2_44_6 ( .A(\ab[44][6] ), .B(\CARRYB[43][6] ), .CI(\SUMB[43][7] ), 
        .CO(\CARRYB[44][6] ), .S(\SUMB[44][6] ) );
  FA1A S2_44_7 ( .A(\ab[44][7] ), .B(\CARRYB[43][7] ), .CI(\SUMB[43][8] ), 
        .CO(\CARRYB[44][7] ), .S(\SUMB[44][7] ) );
  FA1A S2_44_5 ( .A(\ab[44][5] ), .B(\CARRYB[43][5] ), .CI(\SUMB[43][6] ), 
        .CO(\CARRYB[44][5] ), .S(\SUMB[44][5] ) );
  FA1A S2_44_4 ( .A(\ab[44][4] ), .B(\CARRYB[43][4] ), .CI(\SUMB[43][5] ), 
        .CO(\CARRYB[44][4] ), .S(\SUMB[44][4] ) );
  FA1A S2_44_1 ( .A(\ab[44][1] ), .B(\CARRYB[43][1] ), .CI(\SUMB[43][2] ), 
        .CO(\CARRYB[44][1] ), .S(\SUMB[44][1] ) );
  FA1A S2_44_2 ( .A(\ab[44][2] ), .B(\CARRYB[43][2] ), .CI(\SUMB[43][3] ), 
        .CO(\CARRYB[44][2] ), .S(\SUMB[44][2] ) );
  FA1A S2_44_3 ( .A(\ab[44][3] ), .B(\CARRYB[43][3] ), .CI(\SUMB[43][4] ), 
        .CO(\CARRYB[44][3] ), .S(\SUMB[44][3] ) );
  FA1A S2_44_14 ( .A(\ab[44][14] ), .B(\CARRYB[43][14] ), .CI(\SUMB[43][15] ), 
        .CO(\CARRYB[44][14] ), .S(\SUMB[44][14] ) );
  FA1A S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1A S2_41_18 ( .A(\ab[41][18] ), .B(\CARRYB[40][18] ), .CI(\SUMB[40][19] ), 
        .CO(\CARRYB[41][18] ), .S(\SUMB[41][18] ) );
  FA1A S2_41_19 ( .A(\ab[41][19] ), .B(\CARRYB[40][19] ), .CI(\SUMB[40][20] ), 
        .CO(\CARRYB[41][19] ), .S(\SUMB[41][19] ) );
  FA1A S2_43_8 ( .A(\ab[43][8] ), .B(\CARRYB[42][8] ), .CI(\SUMB[42][9] ), 
        .CO(\CARRYB[43][8] ), .S(\SUMB[43][8] ) );
  FA1A S2_43_9 ( .A(\ab[43][9] ), .B(\CARRYB[42][9] ), .CI(\SUMB[42][10] ), 
        .CO(\CARRYB[43][9] ), .S(\SUMB[43][9] ) );
  FA1A S2_43_10 ( .A(\ab[43][10] ), .B(\CARRYB[42][10] ), .CI(\SUMB[42][11] ), 
        .CO(\CARRYB[43][10] ), .S(\SUMB[43][10] ) );
  FA1A S2_43_11 ( .A(\ab[43][11] ), .B(\CARRYB[42][11] ), .CI(\SUMB[42][12] ), 
        .CO(\CARRYB[43][11] ), .S(\SUMB[43][11] ) );
  FA1A S2_43_12 ( .A(\ab[43][12] ), .B(\CARRYB[42][12] ), .CI(\SUMB[42][13] ), 
        .CO(\CARRYB[43][12] ), .S(\SUMB[43][12] ) );
  FA1A S2_43_13 ( .A(\ab[43][13] ), .B(\CARRYB[42][13] ), .CI(\SUMB[42][14] ), 
        .CO(\CARRYB[43][13] ), .S(\SUMB[43][13] ) );
  FA1A S2_43_14 ( .A(\ab[43][14] ), .B(\CARRYB[42][14] ), .CI(\SUMB[42][15] ), 
        .CO(\CARRYB[43][14] ), .S(\SUMB[43][14] ) );
  FA1A S2_43_6 ( .A(\ab[43][6] ), .B(\CARRYB[42][6] ), .CI(\SUMB[42][7] ), 
        .CO(\CARRYB[43][6] ), .S(\SUMB[43][6] ) );
  FA1A S2_43_7 ( .A(\ab[43][7] ), .B(\CARRYB[42][7] ), .CI(\SUMB[42][8] ), 
        .CO(\CARRYB[43][7] ), .S(\SUMB[43][7] ) );
  FA1A S2_43_5 ( .A(\ab[43][5] ), .B(\CARRYB[42][5] ), .CI(\SUMB[42][6] ), 
        .CO(\CARRYB[43][5] ), .S(\SUMB[43][5] ) );
  FA1A S2_43_4 ( .A(\ab[43][4] ), .B(\CARRYB[42][4] ), .CI(\SUMB[42][5] ), 
        .CO(\CARRYB[43][4] ), .S(\SUMB[43][4] ) );
  FA1A S2_43_1 ( .A(\ab[43][1] ), .B(\CARRYB[42][1] ), .CI(\SUMB[42][2] ), 
        .CO(\CARRYB[43][1] ), .S(\SUMB[43][1] ) );
  FA1A S2_43_2 ( .A(\ab[43][2] ), .B(\CARRYB[42][2] ), .CI(\SUMB[42][3] ), 
        .CO(\CARRYB[43][2] ), .S(\SUMB[43][2] ) );
  FA1A S2_43_3 ( .A(\ab[43][3] ), .B(\CARRYB[42][3] ), .CI(\SUMB[42][4] ), 
        .CO(\CARRYB[43][3] ), .S(\SUMB[43][3] ) );
  FA1A S2_43_15 ( .A(\ab[43][15] ), .B(\CARRYB[42][15] ), .CI(\SUMB[42][16] ), 
        .CO(\CARRYB[43][15] ), .S(\SUMB[43][15] ) );
  FA1A S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_40_19 ( .A(\ab[40][19] ), .B(\CARRYB[39][19] ), .CI(\SUMB[39][20] ), 
        .CO(\CARRYB[40][19] ), .S(\SUMB[40][19] ) );
  FA1A S3_40_20 ( .A(\ab[40][20] ), .B(\CARRYB[39][20] ), .CI(\ab[39][21] ), 
        .CO(\CARRYB[40][20] ), .S(\SUMB[40][20] ) );
  FA1A S2_42_8 ( .A(\ab[42][8] ), .B(\CARRYB[41][8] ), .CI(\SUMB[41][9] ), 
        .CO(\CARRYB[42][8] ), .S(\SUMB[42][8] ) );
  FA1A S2_42_9 ( .A(\ab[42][9] ), .B(\CARRYB[41][9] ), .CI(\SUMB[41][10] ), 
        .CO(\CARRYB[42][9] ), .S(\SUMB[42][9] ) );
  FA1A S2_42_10 ( .A(\ab[42][10] ), .B(\CARRYB[41][10] ), .CI(\SUMB[41][11] ), 
        .CO(\CARRYB[42][10] ), .S(\SUMB[42][10] ) );
  FA1A S2_42_11 ( .A(\ab[42][11] ), .B(\CARRYB[41][11] ), .CI(\SUMB[41][12] ), 
        .CO(\CARRYB[42][11] ), .S(\SUMB[42][11] ) );
  FA1A S2_42_12 ( .A(\ab[42][12] ), .B(\CARRYB[41][12] ), .CI(\SUMB[41][13] ), 
        .CO(\CARRYB[42][12] ), .S(\SUMB[42][12] ) );
  FA1A S2_42_13 ( .A(\ab[42][13] ), .B(\CARRYB[41][13] ), .CI(\SUMB[41][14] ), 
        .CO(\CARRYB[42][13] ), .S(\SUMB[42][13] ) );
  FA1A S2_42_14 ( .A(\ab[42][14] ), .B(\CARRYB[41][14] ), .CI(\SUMB[41][15] ), 
        .CO(\CARRYB[42][14] ), .S(\SUMB[42][14] ) );
  FA1A S2_42_15 ( .A(\ab[42][15] ), .B(\CARRYB[41][15] ), .CI(\SUMB[41][16] ), 
        .CO(\CARRYB[42][15] ), .S(\SUMB[42][15] ) );
  FA1A S2_42_6 ( .A(\ab[42][6] ), .B(\CARRYB[41][6] ), .CI(\SUMB[41][7] ), 
        .CO(\CARRYB[42][6] ), .S(\SUMB[42][6] ) );
  FA1A S2_42_7 ( .A(\ab[42][7] ), .B(\CARRYB[41][7] ), .CI(\SUMB[41][8] ), 
        .CO(\CARRYB[42][7] ), .S(\SUMB[42][7] ) );
  FA1A S2_42_5 ( .A(\ab[42][5] ), .B(\CARRYB[41][5] ), .CI(\SUMB[41][6] ), 
        .CO(\CARRYB[42][5] ), .S(\SUMB[42][5] ) );
  FA1A S2_42_4 ( .A(\ab[42][4] ), .B(\CARRYB[41][4] ), .CI(\SUMB[41][5] ), 
        .CO(\CARRYB[42][4] ), .S(\SUMB[42][4] ) );
  FA1A S2_42_1 ( .A(\ab[42][1] ), .B(\CARRYB[41][1] ), .CI(\SUMB[41][2] ), 
        .CO(\CARRYB[42][1] ), .S(\SUMB[42][1] ) );
  FA1A S2_42_2 ( .A(\ab[42][2] ), .B(\CARRYB[41][2] ), .CI(\SUMB[41][3] ), 
        .CO(\CARRYB[42][2] ), .S(\SUMB[42][2] ) );
  FA1A S2_42_3 ( .A(\ab[42][3] ), .B(\CARRYB[41][3] ), .CI(\SUMB[41][4] ), 
        .CO(\CARRYB[42][3] ), .S(\SUMB[42][3] ) );
  FA1A S2_42_16 ( .A(\ab[42][16] ), .B(\CARRYB[41][16] ), .CI(\SUMB[41][17] ), 
        .CO(\CARRYB[42][16] ), .S(\SUMB[42][16] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S3_39_20 ( .A(\ab[39][20] ), .B(\CARRYB[38][20] ), .CI(\ab[38][21] ), 
        .CO(\CARRYB[39][20] ), .S(\SUMB[39][20] ) );
  FA1A S2_41_8 ( .A(\ab[41][8] ), .B(\CARRYB[40][8] ), .CI(\SUMB[40][9] ), 
        .CO(\CARRYB[41][8] ), .S(\SUMB[41][8] ) );
  FA1A S2_41_9 ( .A(\ab[41][9] ), .B(\CARRYB[40][9] ), .CI(\SUMB[40][10] ), 
        .CO(\CARRYB[41][9] ), .S(\SUMB[41][9] ) );
  FA1A S2_41_10 ( .A(\ab[41][10] ), .B(\CARRYB[40][10] ), .CI(\SUMB[40][11] ), 
        .CO(\CARRYB[41][10] ), .S(\SUMB[41][10] ) );
  FA1A S2_41_11 ( .A(\ab[41][11] ), .B(\CARRYB[40][11] ), .CI(\SUMB[40][12] ), 
        .CO(\CARRYB[41][11] ), .S(\SUMB[41][11] ) );
  FA1A S2_41_12 ( .A(\ab[41][12] ), .B(\CARRYB[40][12] ), .CI(\SUMB[40][13] ), 
        .CO(\CARRYB[41][12] ), .S(\SUMB[41][12] ) );
  FA1A S2_41_13 ( .A(\ab[41][13] ), .B(\CARRYB[40][13] ), .CI(\SUMB[40][14] ), 
        .CO(\CARRYB[41][13] ), .S(\SUMB[41][13] ) );
  FA1A S2_41_14 ( .A(\ab[41][14] ), .B(\CARRYB[40][14] ), .CI(\SUMB[40][15] ), 
        .CO(\CARRYB[41][14] ), .S(\SUMB[41][14] ) );
  FA1A S2_41_15 ( .A(\ab[41][15] ), .B(\CARRYB[40][15] ), .CI(\SUMB[40][16] ), 
        .CO(\CARRYB[41][15] ), .S(\SUMB[41][15] ) );
  FA1A S2_41_16 ( .A(\ab[41][16] ), .B(\CARRYB[40][16] ), .CI(\SUMB[40][17] ), 
        .CO(\CARRYB[41][16] ), .S(\SUMB[41][16] ) );
  FA1A S2_41_6 ( .A(\ab[41][6] ), .B(\CARRYB[40][6] ), .CI(\SUMB[40][7] ), 
        .CO(\CARRYB[41][6] ), .S(\SUMB[41][6] ) );
  FA1A S2_41_7 ( .A(\ab[41][7] ), .B(\CARRYB[40][7] ), .CI(\SUMB[40][8] ), 
        .CO(\CARRYB[41][7] ), .S(\SUMB[41][7] ) );
  FA1A S2_41_5 ( .A(\ab[41][5] ), .B(\CARRYB[40][5] ), .CI(\SUMB[40][6] ), 
        .CO(\CARRYB[41][5] ), .S(\SUMB[41][5] ) );
  FA1A S2_41_4 ( .A(\ab[41][4] ), .B(\CARRYB[40][4] ), .CI(\SUMB[40][5] ), 
        .CO(\CARRYB[41][4] ), .S(\SUMB[41][4] ) );
  FA1A S2_41_1 ( .A(\ab[41][1] ), .B(\CARRYB[40][1] ), .CI(\SUMB[40][2] ), 
        .CO(\CARRYB[41][1] ), .S(\SUMB[41][1] ) );
  FA1A S2_41_2 ( .A(\ab[41][2] ), .B(\CARRYB[40][2] ), .CI(\SUMB[40][3] ), 
        .CO(\CARRYB[41][2] ), .S(\SUMB[41][2] ) );
  FA1A S2_41_3 ( .A(\ab[41][3] ), .B(\CARRYB[40][3] ), .CI(\SUMB[40][4] ), 
        .CO(\CARRYB[41][3] ), .S(\SUMB[41][3] ) );
  FA1A S2_41_17 ( .A(\ab[41][17] ), .B(\CARRYB[40][17] ), .CI(\SUMB[40][18] ), 
        .CO(\CARRYB[41][17] ), .S(\SUMB[41][17] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_40_8 ( .A(\ab[40][8] ), .B(\CARRYB[39][8] ), .CI(\SUMB[39][9] ), 
        .CO(\CARRYB[40][8] ), .S(\SUMB[40][8] ) );
  FA1A S2_40_9 ( .A(\ab[40][9] ), .B(\CARRYB[39][9] ), .CI(\SUMB[39][10] ), 
        .CO(\CARRYB[40][9] ), .S(\SUMB[40][9] ) );
  FA1A S2_40_10 ( .A(\ab[40][10] ), .B(\CARRYB[39][10] ), .CI(\SUMB[39][11] ), 
        .CO(\CARRYB[40][10] ), .S(\SUMB[40][10] ) );
  FA1A S2_40_11 ( .A(\ab[40][11] ), .B(\CARRYB[39][11] ), .CI(\SUMB[39][12] ), 
        .CO(\CARRYB[40][11] ), .S(\SUMB[40][11] ) );
  FA1A S2_40_12 ( .A(\ab[40][12] ), .B(\CARRYB[39][12] ), .CI(\SUMB[39][13] ), 
        .CO(\CARRYB[40][12] ), .S(\SUMB[40][12] ) );
  FA1A S2_40_13 ( .A(\ab[40][13] ), .B(\CARRYB[39][13] ), .CI(\SUMB[39][14] ), 
        .CO(\CARRYB[40][13] ), .S(\SUMB[40][13] ) );
  FA1A S2_40_14 ( .A(\ab[40][14] ), .B(\CARRYB[39][14] ), .CI(\SUMB[39][15] ), 
        .CO(\CARRYB[40][14] ), .S(\SUMB[40][14] ) );
  FA1A S2_40_15 ( .A(\ab[40][15] ), .B(\CARRYB[39][15] ), .CI(\SUMB[39][16] ), 
        .CO(\CARRYB[40][15] ), .S(\SUMB[40][15] ) );
  FA1A S2_40_16 ( .A(\ab[40][16] ), .B(\CARRYB[39][16] ), .CI(\SUMB[39][17] ), 
        .CO(\CARRYB[40][16] ), .S(\SUMB[40][16] ) );
  FA1A S2_40_17 ( .A(\ab[40][17] ), .B(\CARRYB[39][17] ), .CI(\SUMB[39][18] ), 
        .CO(\CARRYB[40][17] ), .S(\SUMB[40][17] ) );
  FA1A S2_40_6 ( .A(\ab[40][6] ), .B(\CARRYB[39][6] ), .CI(\SUMB[39][7] ), 
        .CO(\CARRYB[40][6] ), .S(\SUMB[40][6] ) );
  FA1A S2_40_7 ( .A(\ab[40][7] ), .B(\CARRYB[39][7] ), .CI(\SUMB[39][8] ), 
        .CO(\CARRYB[40][7] ), .S(\SUMB[40][7] ) );
  FA1A S2_40_5 ( .A(\ab[40][5] ), .B(\CARRYB[39][5] ), .CI(\SUMB[39][6] ), 
        .CO(\CARRYB[40][5] ), .S(\SUMB[40][5] ) );
  FA1A S2_40_4 ( .A(\ab[40][4] ), .B(\CARRYB[39][4] ), .CI(\SUMB[39][5] ), 
        .CO(\CARRYB[40][4] ), .S(\SUMB[40][4] ) );
  FA1A S2_40_1 ( .A(\ab[40][1] ), .B(\CARRYB[39][1] ), .CI(\SUMB[39][2] ), 
        .CO(\CARRYB[40][1] ), .S(\SUMB[40][1] ) );
  FA1A S2_40_2 ( .A(\ab[40][2] ), .B(\CARRYB[39][2] ), .CI(\SUMB[39][3] ), 
        .CO(\CARRYB[40][2] ), .S(\SUMB[40][2] ) );
  FA1A S2_40_3 ( .A(\ab[40][3] ), .B(\CARRYB[39][3] ), .CI(\SUMB[39][4] ), 
        .CO(\CARRYB[40][3] ), .S(\SUMB[40][3] ) );
  FA1A S2_40_18 ( .A(\ab[40][18] ), .B(\CARRYB[39][18] ), .CI(\SUMB[39][19] ), 
        .CO(\CARRYB[40][18] ), .S(\SUMB[40][18] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_39_8 ( .A(\ab[39][8] ), .B(\CARRYB[38][8] ), .CI(\SUMB[38][9] ), 
        .CO(\CARRYB[39][8] ), .S(\SUMB[39][8] ) );
  FA1A S2_39_9 ( .A(\ab[39][9] ), .B(\CARRYB[38][9] ), .CI(\SUMB[38][10] ), 
        .CO(\CARRYB[39][9] ), .S(\SUMB[39][9] ) );
  FA1A S2_39_10 ( .A(\ab[39][10] ), .B(\CARRYB[38][10] ), .CI(\SUMB[38][11] ), 
        .CO(\CARRYB[39][10] ), .S(\SUMB[39][10] ) );
  FA1A S2_39_11 ( .A(\ab[39][11] ), .B(\CARRYB[38][11] ), .CI(\SUMB[38][12] ), 
        .CO(\CARRYB[39][11] ), .S(\SUMB[39][11] ) );
  FA1A S2_39_12 ( .A(\ab[39][12] ), .B(\CARRYB[38][12] ), .CI(\SUMB[38][13] ), 
        .CO(\CARRYB[39][12] ), .S(\SUMB[39][12] ) );
  FA1A S2_39_13 ( .A(\ab[39][13] ), .B(\CARRYB[38][13] ), .CI(\SUMB[38][14] ), 
        .CO(\CARRYB[39][13] ), .S(\SUMB[39][13] ) );
  FA1A S2_39_14 ( .A(\ab[39][14] ), .B(\CARRYB[38][14] ), .CI(\SUMB[38][15] ), 
        .CO(\CARRYB[39][14] ), .S(\SUMB[39][14] ) );
  FA1A S2_39_15 ( .A(\ab[39][15] ), .B(\CARRYB[38][15] ), .CI(\SUMB[38][16] ), 
        .CO(\CARRYB[39][15] ), .S(\SUMB[39][15] ) );
  FA1A S2_39_16 ( .A(\ab[39][16] ), .B(\CARRYB[38][16] ), .CI(\SUMB[38][17] ), 
        .CO(\CARRYB[39][16] ), .S(\SUMB[39][16] ) );
  FA1A S2_39_17 ( .A(\ab[39][17] ), .B(\CARRYB[38][17] ), .CI(\SUMB[38][18] ), 
        .CO(\CARRYB[39][17] ), .S(\SUMB[39][17] ) );
  FA1A S2_39_18 ( .A(\ab[39][18] ), .B(\CARRYB[38][18] ), .CI(\SUMB[38][19] ), 
        .CO(\CARRYB[39][18] ), .S(\SUMB[39][18] ) );
  FA1A S2_39_6 ( .A(\ab[39][6] ), .B(\CARRYB[38][6] ), .CI(\SUMB[38][7] ), 
        .CO(\CARRYB[39][6] ), .S(\SUMB[39][6] ) );
  FA1A S2_39_7 ( .A(\ab[39][7] ), .B(\CARRYB[38][7] ), .CI(\SUMB[38][8] ), 
        .CO(\CARRYB[39][7] ), .S(\SUMB[39][7] ) );
  FA1A S2_39_5 ( .A(\ab[39][5] ), .B(\CARRYB[38][5] ), .CI(\SUMB[38][6] ), 
        .CO(\CARRYB[39][5] ), .S(\SUMB[39][5] ) );
  FA1A S2_39_4 ( .A(\ab[39][4] ), .B(\CARRYB[38][4] ), .CI(\SUMB[38][5] ), 
        .CO(\CARRYB[39][4] ), .S(\SUMB[39][4] ) );
  FA1A S2_39_1 ( .A(\ab[39][1] ), .B(\CARRYB[38][1] ), .CI(\SUMB[38][2] ), 
        .CO(\CARRYB[39][1] ), .S(\SUMB[39][1] ) );
  FA1A S2_39_2 ( .A(\ab[39][2] ), .B(\CARRYB[38][2] ), .CI(\SUMB[38][3] ), 
        .CO(\CARRYB[39][2] ), .S(\SUMB[39][2] ) );
  FA1A S2_39_3 ( .A(\ab[39][3] ), .B(\CARRYB[38][3] ), .CI(\SUMB[38][4] ), 
        .CO(\CARRYB[39][3] ), .S(\SUMB[39][3] ) );
  FA1A S2_39_19 ( .A(\ab[39][19] ), .B(\CARRYB[38][19] ), .CI(\SUMB[38][20] ), 
        .CO(\CARRYB[39][19] ), .S(\SUMB[39][19] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_38_8 ( .A(\ab[38][8] ), .B(\CARRYB[37][8] ), .CI(\SUMB[37][9] ), 
        .CO(\CARRYB[38][8] ), .S(\SUMB[38][8] ) );
  FA1A S2_38_9 ( .A(\ab[38][9] ), .B(\CARRYB[37][9] ), .CI(\SUMB[37][10] ), 
        .CO(\CARRYB[38][9] ), .S(\SUMB[38][9] ) );
  FA1A S2_38_10 ( .A(\ab[38][10] ), .B(\CARRYB[37][10] ), .CI(\SUMB[37][11] ), 
        .CO(\CARRYB[38][10] ), .S(\SUMB[38][10] ) );
  FA1A S2_38_11 ( .A(\ab[38][11] ), .B(\CARRYB[37][11] ), .CI(\SUMB[37][12] ), 
        .CO(\CARRYB[38][11] ), .S(\SUMB[38][11] ) );
  FA1A S2_38_12 ( .A(\ab[38][12] ), .B(\CARRYB[37][12] ), .CI(\SUMB[37][13] ), 
        .CO(\CARRYB[38][12] ), .S(\SUMB[38][12] ) );
  FA1A S2_38_13 ( .A(\ab[38][13] ), .B(\CARRYB[37][13] ), .CI(\SUMB[37][14] ), 
        .CO(\CARRYB[38][13] ), .S(\SUMB[38][13] ) );
  FA1A S2_38_14 ( .A(\ab[38][14] ), .B(\CARRYB[37][14] ), .CI(\SUMB[37][15] ), 
        .CO(\CARRYB[38][14] ), .S(\SUMB[38][14] ) );
  FA1A S2_38_15 ( .A(\ab[38][15] ), .B(\CARRYB[37][15] ), .CI(\SUMB[37][16] ), 
        .CO(\CARRYB[38][15] ), .S(\SUMB[38][15] ) );
  FA1A S2_38_16 ( .A(\ab[38][16] ), .B(\CARRYB[37][16] ), .CI(\SUMB[37][17] ), 
        .CO(\CARRYB[38][16] ), .S(\SUMB[38][16] ) );
  FA1A S2_38_17 ( .A(\ab[38][17] ), .B(\CARRYB[37][17] ), .CI(\SUMB[37][18] ), 
        .CO(\CARRYB[38][17] ), .S(\SUMB[38][17] ) );
  FA1A S2_38_18 ( .A(\ab[38][18] ), .B(\CARRYB[37][18] ), .CI(\SUMB[37][19] ), 
        .CO(\CARRYB[38][18] ), .S(\SUMB[38][18] ) );
  FA1A S2_38_19 ( .A(\ab[38][19] ), .B(\CARRYB[37][19] ), .CI(\SUMB[37][20] ), 
        .CO(\CARRYB[38][19] ), .S(\SUMB[38][19] ) );
  FA1A S2_38_6 ( .A(\ab[38][6] ), .B(\CARRYB[37][6] ), .CI(\SUMB[37][7] ), 
        .CO(\CARRYB[38][6] ), .S(\SUMB[38][6] ) );
  FA1A S2_38_7 ( .A(\ab[38][7] ), .B(\CARRYB[37][7] ), .CI(\SUMB[37][8] ), 
        .CO(\CARRYB[38][7] ), .S(\SUMB[38][7] ) );
  FA1A S2_38_5 ( .A(\ab[38][5] ), .B(\CARRYB[37][5] ), .CI(\SUMB[37][6] ), 
        .CO(\CARRYB[38][5] ), .S(\SUMB[38][5] ) );
  FA1A S2_38_4 ( .A(\ab[38][4] ), .B(\CARRYB[37][4] ), .CI(\SUMB[37][5] ), 
        .CO(\CARRYB[38][4] ), .S(\SUMB[38][4] ) );
  FA1A S2_38_1 ( .A(\ab[38][1] ), .B(\CARRYB[37][1] ), .CI(\SUMB[37][2] ), 
        .CO(\CARRYB[38][1] ), .S(\SUMB[38][1] ) );
  FA1A S2_38_2 ( .A(\ab[38][2] ), .B(\CARRYB[37][2] ), .CI(\SUMB[37][3] ), 
        .CO(\CARRYB[38][2] ), .S(\SUMB[38][2] ) );
  FA1A S2_38_3 ( .A(\ab[38][3] ), .B(\CARRYB[37][3] ), .CI(\SUMB[37][4] ), 
        .CO(\CARRYB[38][3] ), .S(\SUMB[38][3] ) );
  FA1A S3_38_20 ( .A(\ab[38][20] ), .B(\CARRYB[37][20] ), .CI(\ab[37][21] ), 
        .CO(\CARRYB[38][20] ), .S(\SUMB[38][20] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_37_8 ( .A(\ab[37][8] ), .B(\CARRYB[36][8] ), .CI(\SUMB[36][9] ), 
        .CO(\CARRYB[37][8] ), .S(\SUMB[37][8] ) );
  FA1A S2_37_9 ( .A(\ab[37][9] ), .B(\CARRYB[36][9] ), .CI(\SUMB[36][10] ), 
        .CO(\CARRYB[37][9] ), .S(\SUMB[37][9] ) );
  FA1A S2_37_10 ( .A(\ab[37][10] ), .B(\CARRYB[36][10] ), .CI(\SUMB[36][11] ), 
        .CO(\CARRYB[37][10] ), .S(\SUMB[37][10] ) );
  FA1A S2_37_11 ( .A(\ab[37][11] ), .B(\CARRYB[36][11] ), .CI(\SUMB[36][12] ), 
        .CO(\CARRYB[37][11] ), .S(\SUMB[37][11] ) );
  FA1A S2_37_12 ( .A(\ab[37][12] ), .B(\CARRYB[36][12] ), .CI(\SUMB[36][13] ), 
        .CO(\CARRYB[37][12] ), .S(\SUMB[37][12] ) );
  FA1A S2_37_13 ( .A(\ab[37][13] ), .B(\CARRYB[36][13] ), .CI(\SUMB[36][14] ), 
        .CO(\CARRYB[37][13] ), .S(\SUMB[37][13] ) );
  FA1A S2_37_14 ( .A(\ab[37][14] ), .B(\CARRYB[36][14] ), .CI(\SUMB[36][15] ), 
        .CO(\CARRYB[37][14] ), .S(\SUMB[37][14] ) );
  FA1A S2_37_15 ( .A(\ab[37][15] ), .B(\CARRYB[36][15] ), .CI(\SUMB[36][16] ), 
        .CO(\CARRYB[37][15] ), .S(\SUMB[37][15] ) );
  FA1A S2_37_16 ( .A(\ab[37][16] ), .B(\CARRYB[36][16] ), .CI(\SUMB[36][17] ), 
        .CO(\CARRYB[37][16] ), .S(\SUMB[37][16] ) );
  FA1A S2_37_17 ( .A(\ab[37][17] ), .B(\CARRYB[36][17] ), .CI(\SUMB[36][18] ), 
        .CO(\CARRYB[37][17] ), .S(\SUMB[37][17] ) );
  FA1A S2_37_18 ( .A(\ab[37][18] ), .B(\CARRYB[36][18] ), .CI(\SUMB[36][19] ), 
        .CO(\CARRYB[37][18] ), .S(\SUMB[37][18] ) );
  FA1A S2_37_19 ( .A(\ab[37][19] ), .B(\CARRYB[36][19] ), .CI(\SUMB[36][20] ), 
        .CO(\CARRYB[37][19] ), .S(\SUMB[37][19] ) );
  FA1A S3_37_20 ( .A(\ab[37][20] ), .B(\CARRYB[36][20] ), .CI(\ab[36][21] ), 
        .CO(\CARRYB[37][20] ), .S(\SUMB[37][20] ) );
  FA1A S2_37_6 ( .A(\ab[37][6] ), .B(\CARRYB[36][6] ), .CI(\SUMB[36][7] ), 
        .CO(\CARRYB[37][6] ), .S(\SUMB[37][6] ) );
  FA1A S2_37_7 ( .A(\ab[37][7] ), .B(\CARRYB[36][7] ), .CI(\SUMB[36][8] ), 
        .CO(\CARRYB[37][7] ), .S(\SUMB[37][7] ) );
  FA1A S2_37_5 ( .A(\ab[37][5] ), .B(\CARRYB[36][5] ), .CI(\SUMB[36][6] ), 
        .CO(\CARRYB[37][5] ), .S(\SUMB[37][5] ) );
  FA1A S2_37_4 ( .A(\ab[37][4] ), .B(\CARRYB[36][4] ), .CI(\SUMB[36][5] ), 
        .CO(\CARRYB[37][4] ), .S(\SUMB[37][4] ) );
  FA1A S2_37_1 ( .A(\ab[37][1] ), .B(\CARRYB[36][1] ), .CI(\SUMB[36][2] ), 
        .CO(\CARRYB[37][1] ), .S(\SUMB[37][1] ) );
  FA1A S2_37_2 ( .A(\ab[37][2] ), .B(\CARRYB[36][2] ), .CI(\SUMB[36][3] ), 
        .CO(\CARRYB[37][2] ), .S(\SUMB[37][2] ) );
  FA1A S2_37_3 ( .A(\ab[37][3] ), .B(\CARRYB[36][3] ), .CI(\SUMB[36][4] ), 
        .CO(\CARRYB[37][3] ), .S(\SUMB[37][3] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_36_8 ( .A(\ab[36][8] ), .B(\CARRYB[35][8] ), .CI(\SUMB[35][9] ), 
        .CO(\CARRYB[36][8] ), .S(\SUMB[36][8] ) );
  FA1A S2_36_9 ( .A(\ab[36][9] ), .B(\CARRYB[35][9] ), .CI(\SUMB[35][10] ), 
        .CO(\CARRYB[36][9] ), .S(\SUMB[36][9] ) );
  FA1A S2_36_10 ( .A(\ab[36][10] ), .B(\CARRYB[35][10] ), .CI(\SUMB[35][11] ), 
        .CO(\CARRYB[36][10] ), .S(\SUMB[36][10] ) );
  FA1A S2_36_11 ( .A(\ab[36][11] ), .B(\CARRYB[35][11] ), .CI(\SUMB[35][12] ), 
        .CO(\CARRYB[36][11] ), .S(\SUMB[36][11] ) );
  FA1A S2_36_12 ( .A(\ab[36][12] ), .B(\CARRYB[35][12] ), .CI(\SUMB[35][13] ), 
        .CO(\CARRYB[36][12] ), .S(\SUMB[36][12] ) );
  FA1A S2_36_13 ( .A(\ab[36][13] ), .B(\CARRYB[35][13] ), .CI(\SUMB[35][14] ), 
        .CO(\CARRYB[36][13] ), .S(\SUMB[36][13] ) );
  FA1A S2_36_14 ( .A(\ab[36][14] ), .B(\CARRYB[35][14] ), .CI(\SUMB[35][15] ), 
        .CO(\CARRYB[36][14] ), .S(\SUMB[36][14] ) );
  FA1A S2_36_15 ( .A(\ab[36][15] ), .B(\CARRYB[35][15] ), .CI(\SUMB[35][16] ), 
        .CO(\CARRYB[36][15] ), .S(\SUMB[36][15] ) );
  FA1A S2_36_16 ( .A(\ab[36][16] ), .B(\CARRYB[35][16] ), .CI(\SUMB[35][17] ), 
        .CO(\CARRYB[36][16] ), .S(\SUMB[36][16] ) );
  FA1A S2_36_17 ( .A(\ab[36][17] ), .B(\CARRYB[35][17] ), .CI(\SUMB[35][18] ), 
        .CO(\CARRYB[36][17] ), .S(\SUMB[36][17] ) );
  FA1A S2_36_18 ( .A(\ab[36][18] ), .B(\CARRYB[35][18] ), .CI(\SUMB[35][19] ), 
        .CO(\CARRYB[36][18] ), .S(\SUMB[36][18] ) );
  FA1A S2_36_19 ( .A(\ab[36][19] ), .B(\CARRYB[35][19] ), .CI(\SUMB[35][20] ), 
        .CO(\CARRYB[36][19] ), .S(\SUMB[36][19] ) );
  FA1A S3_36_20 ( .A(\ab[36][20] ), .B(\CARRYB[35][20] ), .CI(\ab[35][21] ), 
        .CO(\CARRYB[36][20] ), .S(\SUMB[36][20] ) );
  FA1A S2_36_6 ( .A(\ab[36][6] ), .B(\CARRYB[35][6] ), .CI(\SUMB[35][7] ), 
        .CO(\CARRYB[36][6] ), .S(\SUMB[36][6] ) );
  FA1A S2_36_7 ( .A(\ab[36][7] ), .B(\CARRYB[35][7] ), .CI(\SUMB[35][8] ), 
        .CO(\CARRYB[36][7] ), .S(\SUMB[36][7] ) );
  FA1A S2_36_5 ( .A(\ab[36][5] ), .B(\CARRYB[35][5] ), .CI(\SUMB[35][6] ), 
        .CO(\CARRYB[36][5] ), .S(\SUMB[36][5] ) );
  FA1A S2_36_4 ( .A(\ab[36][4] ), .B(\CARRYB[35][4] ), .CI(\SUMB[35][5] ), 
        .CO(\CARRYB[36][4] ), .S(\SUMB[36][4] ) );
  FA1A S2_36_2 ( .A(\ab[36][2] ), .B(\CARRYB[35][2] ), .CI(\SUMB[35][3] ), 
        .CO(\CARRYB[36][2] ), .S(\SUMB[36][2] ) );
  FA1A S2_36_3 ( .A(\ab[36][3] ), .B(\CARRYB[35][3] ), .CI(\SUMB[35][4] ), 
        .CO(\CARRYB[36][3] ), .S(\SUMB[36][3] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_35_8 ( .A(\ab[35][8] ), .B(\CARRYB[34][8] ), .CI(\SUMB[34][9] ), 
        .CO(\CARRYB[35][8] ), .S(\SUMB[35][8] ) );
  FA1A S2_35_9 ( .A(\ab[35][9] ), .B(\CARRYB[34][9] ), .CI(\SUMB[34][10] ), 
        .CO(\CARRYB[35][9] ), .S(\SUMB[35][9] ) );
  FA1A S2_35_10 ( .A(\ab[35][10] ), .B(\CARRYB[34][10] ), .CI(\SUMB[34][11] ), 
        .CO(\CARRYB[35][10] ), .S(\SUMB[35][10] ) );
  FA1A S2_35_11 ( .A(\ab[35][11] ), .B(\CARRYB[34][11] ), .CI(\SUMB[34][12] ), 
        .CO(\CARRYB[35][11] ), .S(\SUMB[35][11] ) );
  FA1A S2_35_12 ( .A(\ab[35][12] ), .B(\CARRYB[34][12] ), .CI(\SUMB[34][13] ), 
        .CO(\CARRYB[35][12] ), .S(\SUMB[35][12] ) );
  FA1A S2_35_13 ( .A(\ab[35][13] ), .B(\CARRYB[34][13] ), .CI(\SUMB[34][14] ), 
        .CO(\CARRYB[35][13] ), .S(\SUMB[35][13] ) );
  FA1A S2_35_14 ( .A(\ab[35][14] ), .B(\CARRYB[34][14] ), .CI(\SUMB[34][15] ), 
        .CO(\CARRYB[35][14] ), .S(\SUMB[35][14] ) );
  FA1A S2_35_15 ( .A(\ab[35][15] ), .B(\CARRYB[34][15] ), .CI(\SUMB[34][16] ), 
        .CO(\CARRYB[35][15] ), .S(\SUMB[35][15] ) );
  FA1A S2_35_16 ( .A(\ab[35][16] ), .B(\CARRYB[34][16] ), .CI(\SUMB[34][17] ), 
        .CO(\CARRYB[35][16] ), .S(\SUMB[35][16] ) );
  FA1A S2_35_17 ( .A(\ab[35][17] ), .B(\CARRYB[34][17] ), .CI(\SUMB[34][18] ), 
        .CO(\CARRYB[35][17] ), .S(\SUMB[35][17] ) );
  FA1A S2_35_18 ( .A(\ab[35][18] ), .B(\CARRYB[34][18] ), .CI(\SUMB[34][19] ), 
        .CO(\CARRYB[35][18] ), .S(\SUMB[35][18] ) );
  FA1A S2_35_19 ( .A(\ab[35][19] ), .B(\CARRYB[34][19] ), .CI(\SUMB[34][20] ), 
        .CO(\CARRYB[35][19] ), .S(\SUMB[35][19] ) );
  FA1A S3_35_20 ( .A(\ab[35][20] ), .B(\CARRYB[34][20] ), .CI(\ab[34][21] ), 
        .CO(\CARRYB[35][20] ), .S(\SUMB[35][20] ) );
  FA1A S2_35_6 ( .A(\ab[35][6] ), .B(\CARRYB[34][6] ), .CI(\SUMB[34][7] ), 
        .CO(\CARRYB[35][6] ), .S(\SUMB[35][6] ) );
  FA1A S2_35_7 ( .A(\ab[35][7] ), .B(\CARRYB[34][7] ), .CI(\SUMB[34][8] ), 
        .CO(\CARRYB[35][7] ), .S(\SUMB[35][7] ) );
  FA1A S2_35_5 ( .A(\ab[35][5] ), .B(\CARRYB[34][5] ), .CI(\SUMB[34][6] ), 
        .CO(\CARRYB[35][5] ), .S(\SUMB[35][5] ) );
  FA1A S2_35_4 ( .A(\ab[35][4] ), .B(\CARRYB[34][4] ), .CI(\SUMB[34][5] ), 
        .CO(\CARRYB[35][4] ), .S(\SUMB[35][4] ) );
  FA1A S2_35_2 ( .A(\ab[35][2] ), .B(\CARRYB[34][2] ), .CI(\SUMB[34][3] ), 
        .CO(\CARRYB[35][2] ), .S(\SUMB[35][2] ) );
  FA1A S2_35_3 ( .A(\ab[35][3] ), .B(\CARRYB[34][3] ), .CI(\SUMB[34][4] ), 
        .CO(\CARRYB[35][3] ), .S(\SUMB[35][3] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_34_8 ( .A(\ab[34][8] ), .B(\CARRYB[33][8] ), .CI(\SUMB[33][9] ), 
        .CO(\CARRYB[34][8] ), .S(\SUMB[34][8] ) );
  FA1A S2_34_9 ( .A(\ab[34][9] ), .B(\CARRYB[33][9] ), .CI(\SUMB[33][10] ), 
        .CO(\CARRYB[34][9] ), .S(\SUMB[34][9] ) );
  FA1A S2_34_10 ( .A(\ab[34][10] ), .B(\CARRYB[33][10] ), .CI(\SUMB[33][11] ), 
        .CO(\CARRYB[34][10] ), .S(\SUMB[34][10] ) );
  FA1A S2_34_11 ( .A(\ab[34][11] ), .B(\CARRYB[33][11] ), .CI(\SUMB[33][12] ), 
        .CO(\CARRYB[34][11] ), .S(\SUMB[34][11] ) );
  FA1A S2_34_12 ( .A(\ab[34][12] ), .B(\CARRYB[33][12] ), .CI(\SUMB[33][13] ), 
        .CO(\CARRYB[34][12] ), .S(\SUMB[34][12] ) );
  FA1A S2_34_13 ( .A(\ab[34][13] ), .B(\CARRYB[33][13] ), .CI(\SUMB[33][14] ), 
        .CO(\CARRYB[34][13] ), .S(\SUMB[34][13] ) );
  FA1A S2_34_14 ( .A(\ab[34][14] ), .B(\CARRYB[33][14] ), .CI(\SUMB[33][15] ), 
        .CO(\CARRYB[34][14] ), .S(\SUMB[34][14] ) );
  FA1A S2_34_15 ( .A(\ab[34][15] ), .B(\CARRYB[33][15] ), .CI(\SUMB[33][16] ), 
        .CO(\CARRYB[34][15] ), .S(\SUMB[34][15] ) );
  FA1A S2_34_16 ( .A(\ab[34][16] ), .B(\CARRYB[33][16] ), .CI(\SUMB[33][17] ), 
        .CO(\CARRYB[34][16] ), .S(\SUMB[34][16] ) );
  FA1A S2_34_17 ( .A(\ab[34][17] ), .B(\CARRYB[33][17] ), .CI(\SUMB[33][18] ), 
        .CO(\CARRYB[34][17] ), .S(\SUMB[34][17] ) );
  FA1A S2_34_18 ( .A(\ab[34][18] ), .B(\CARRYB[33][18] ), .CI(\SUMB[33][19] ), 
        .CO(\CARRYB[34][18] ), .S(\SUMB[34][18] ) );
  FA1A S2_34_19 ( .A(\ab[34][19] ), .B(\CARRYB[33][19] ), .CI(\SUMB[33][20] ), 
        .CO(\CARRYB[34][19] ), .S(\SUMB[34][19] ) );
  FA1A S3_34_20 ( .A(\ab[34][20] ), .B(\CARRYB[33][20] ), .CI(\ab[33][21] ), 
        .CO(\CARRYB[34][20] ), .S(\SUMB[34][20] ) );
  FA1A S2_34_6 ( .A(\ab[34][6] ), .B(\CARRYB[33][6] ), .CI(\SUMB[33][7] ), 
        .CO(\CARRYB[34][6] ), .S(\SUMB[34][6] ) );
  FA1A S2_34_7 ( .A(\ab[34][7] ), .B(\CARRYB[33][7] ), .CI(\SUMB[33][8] ), 
        .CO(\CARRYB[34][7] ), .S(\SUMB[34][7] ) );
  FA1A S2_34_5 ( .A(\ab[34][5] ), .B(\CARRYB[33][5] ), .CI(\SUMB[33][6] ), 
        .CO(\CARRYB[34][5] ), .S(\SUMB[34][5] ) );
  FA1A S2_34_4 ( .A(\ab[34][4] ), .B(\CARRYB[33][4] ), .CI(\SUMB[33][5] ), 
        .CO(\CARRYB[34][4] ), .S(\SUMB[34][4] ) );
  FA1A S2_34_2 ( .A(\ab[34][2] ), .B(\CARRYB[33][2] ), .CI(\SUMB[33][3] ), 
        .CO(\CARRYB[34][2] ), .S(\SUMB[34][2] ) );
  FA1A S2_34_3 ( .A(\ab[34][3] ), .B(\CARRYB[33][3] ), .CI(\SUMB[33][4] ), 
        .CO(\CARRYB[34][3] ), .S(\SUMB[34][3] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_33_8 ( .A(\ab[33][8] ), .B(\CARRYB[32][8] ), .CI(\SUMB[32][9] ), 
        .CO(\CARRYB[33][8] ), .S(\SUMB[33][8] ) );
  FA1A S2_33_9 ( .A(\ab[33][9] ), .B(\CARRYB[32][9] ), .CI(\SUMB[32][10] ), 
        .CO(\CARRYB[33][9] ), .S(\SUMB[33][9] ) );
  FA1A S2_33_10 ( .A(\ab[33][10] ), .B(\CARRYB[32][10] ), .CI(\SUMB[32][11] ), 
        .CO(\CARRYB[33][10] ), .S(\SUMB[33][10] ) );
  FA1A S2_33_11 ( .A(\ab[33][11] ), .B(\CARRYB[32][11] ), .CI(\SUMB[32][12] ), 
        .CO(\CARRYB[33][11] ), .S(\SUMB[33][11] ) );
  FA1A S2_33_12 ( .A(\ab[33][12] ), .B(\CARRYB[32][12] ), .CI(\SUMB[32][13] ), 
        .CO(\CARRYB[33][12] ), .S(\SUMB[33][12] ) );
  FA1A S2_33_13 ( .A(\ab[33][13] ), .B(\CARRYB[32][13] ), .CI(\SUMB[32][14] ), 
        .CO(\CARRYB[33][13] ), .S(\SUMB[33][13] ) );
  FA1A S2_33_14 ( .A(\ab[33][14] ), .B(\CARRYB[32][14] ), .CI(\SUMB[32][15] ), 
        .CO(\CARRYB[33][14] ), .S(\SUMB[33][14] ) );
  FA1A S2_33_15 ( .A(\ab[33][15] ), .B(\CARRYB[32][15] ), .CI(\SUMB[32][16] ), 
        .CO(\CARRYB[33][15] ), .S(\SUMB[33][15] ) );
  FA1A S2_33_16 ( .A(\ab[33][16] ), .B(\CARRYB[32][16] ), .CI(\SUMB[32][17] ), 
        .CO(\CARRYB[33][16] ), .S(\SUMB[33][16] ) );
  FA1A S2_33_17 ( .A(\ab[33][17] ), .B(\CARRYB[32][17] ), .CI(\SUMB[32][18] ), 
        .CO(\CARRYB[33][17] ), .S(\SUMB[33][17] ) );
  FA1A S2_33_18 ( .A(\ab[33][18] ), .B(\CARRYB[32][18] ), .CI(\SUMB[32][19] ), 
        .CO(\CARRYB[33][18] ), .S(\SUMB[33][18] ) );
  FA1A S2_33_19 ( .A(\ab[33][19] ), .B(\CARRYB[32][19] ), .CI(\SUMB[32][20] ), 
        .CO(\CARRYB[33][19] ), .S(\SUMB[33][19] ) );
  FA1A S3_33_20 ( .A(\ab[33][20] ), .B(\CARRYB[32][20] ), .CI(\ab[32][21] ), 
        .CO(\CARRYB[33][20] ), .S(\SUMB[33][20] ) );
  FA1A S2_33_6 ( .A(\ab[33][6] ), .B(\CARRYB[32][6] ), .CI(\SUMB[32][7] ), 
        .CO(\CARRYB[33][6] ), .S(\SUMB[33][6] ) );
  FA1A S2_33_7 ( .A(\ab[33][7] ), .B(\CARRYB[32][7] ), .CI(\SUMB[32][8] ), 
        .CO(\CARRYB[33][7] ), .S(\SUMB[33][7] ) );
  FA1A S2_33_5 ( .A(\ab[33][5] ), .B(\CARRYB[32][5] ), .CI(\SUMB[32][6] ), 
        .CO(\CARRYB[33][5] ), .S(\SUMB[33][5] ) );
  FA1A S2_33_4 ( .A(\ab[33][4] ), .B(\CARRYB[32][4] ), .CI(\SUMB[32][5] ), 
        .CO(\CARRYB[33][4] ), .S(\SUMB[33][4] ) );
  FA1A S2_33_2 ( .A(\ab[33][2] ), .B(\CARRYB[32][2] ), .CI(\SUMB[32][3] ), 
        .CO(\CARRYB[33][2] ), .S(\SUMB[33][2] ) );
  FA1A S2_33_3 ( .A(\ab[33][3] ), .B(\CARRYB[32][3] ), .CI(\SUMB[32][4] ), 
        .CO(\CARRYB[33][3] ), .S(\SUMB[33][3] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_32_8 ( .A(\ab[32][8] ), .B(\CARRYB[31][8] ), .CI(\SUMB[31][9] ), 
        .CO(\CARRYB[32][8] ), .S(\SUMB[32][8] ) );
  FA1A S2_32_9 ( .A(\ab[32][9] ), .B(\CARRYB[31][9] ), .CI(\SUMB[31][10] ), 
        .CO(\CARRYB[32][9] ), .S(\SUMB[32][9] ) );
  FA1A S2_32_10 ( .A(\ab[32][10] ), .B(\CARRYB[31][10] ), .CI(\SUMB[31][11] ), 
        .CO(\CARRYB[32][10] ), .S(\SUMB[32][10] ) );
  FA1A S2_32_11 ( .A(\ab[32][11] ), .B(\CARRYB[31][11] ), .CI(\SUMB[31][12] ), 
        .CO(\CARRYB[32][11] ), .S(\SUMB[32][11] ) );
  FA1A S2_32_12 ( .A(\ab[32][12] ), .B(\CARRYB[31][12] ), .CI(\SUMB[31][13] ), 
        .CO(\CARRYB[32][12] ), .S(\SUMB[32][12] ) );
  FA1A S2_32_13 ( .A(\ab[32][13] ), .B(\CARRYB[31][13] ), .CI(\SUMB[31][14] ), 
        .CO(\CARRYB[32][13] ), .S(\SUMB[32][13] ) );
  FA1A S2_32_14 ( .A(\ab[32][14] ), .B(\CARRYB[31][14] ), .CI(\SUMB[31][15] ), 
        .CO(\CARRYB[32][14] ), .S(\SUMB[32][14] ) );
  FA1A S2_32_15 ( .A(\ab[32][15] ), .B(\CARRYB[31][15] ), .CI(\SUMB[31][16] ), 
        .CO(\CARRYB[32][15] ), .S(\SUMB[32][15] ) );
  FA1A S2_32_16 ( .A(\ab[32][16] ), .B(\CARRYB[31][16] ), .CI(\SUMB[31][17] ), 
        .CO(\CARRYB[32][16] ), .S(\SUMB[32][16] ) );
  FA1A S2_32_17 ( .A(\ab[32][17] ), .B(\CARRYB[31][17] ), .CI(\SUMB[31][18] ), 
        .CO(\CARRYB[32][17] ), .S(\SUMB[32][17] ) );
  FA1A S2_32_18 ( .A(\ab[32][18] ), .B(\CARRYB[31][18] ), .CI(\SUMB[31][19] ), 
        .CO(\CARRYB[32][18] ), .S(\SUMB[32][18] ) );
  FA1A S2_32_19 ( .A(\ab[32][19] ), .B(\CARRYB[31][19] ), .CI(\SUMB[31][20] ), 
        .CO(\CARRYB[32][19] ), .S(\SUMB[32][19] ) );
  FA1A S3_32_20 ( .A(\ab[32][20] ), .B(\CARRYB[31][20] ), .CI(\ab[31][21] ), 
        .CO(\CARRYB[32][20] ), .S(\SUMB[32][20] ) );
  FA1A S2_32_6 ( .A(\ab[32][6] ), .B(\CARRYB[31][6] ), .CI(\SUMB[31][7] ), 
        .CO(\CARRYB[32][6] ), .S(\SUMB[32][6] ) );
  FA1A S2_32_7 ( .A(\ab[32][7] ), .B(\CARRYB[31][7] ), .CI(\SUMB[31][8] ), 
        .CO(\CARRYB[32][7] ), .S(\SUMB[32][7] ) );
  FA1A S2_32_5 ( .A(\ab[32][5] ), .B(\CARRYB[31][5] ), .CI(\SUMB[31][6] ), 
        .CO(\CARRYB[32][5] ), .S(\SUMB[32][5] ) );
  FA1A S2_32_4 ( .A(\ab[32][4] ), .B(\CARRYB[31][4] ), .CI(\SUMB[31][5] ), 
        .CO(\CARRYB[32][4] ), .S(\SUMB[32][4] ) );
  FA1A S2_32_2 ( .A(\ab[32][2] ), .B(\CARRYB[31][2] ), .CI(\SUMB[31][3] ), 
        .CO(\CARRYB[32][2] ), .S(\SUMB[32][2] ) );
  FA1A S2_32_3 ( .A(\ab[32][3] ), .B(\CARRYB[31][3] ), .CI(\SUMB[31][4] ), 
        .CO(\CARRYB[32][3] ), .S(\SUMB[32][3] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_31_8 ( .A(\ab[31][8] ), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), 
        .CO(\CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA1A S2_31_9 ( .A(\ab[31][9] ), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), 
        .CO(\CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA1A S2_31_10 ( .A(\ab[31][10] ), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), 
        .CO(\CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA1A S2_31_11 ( .A(\ab[31][11] ), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), 
        .CO(\CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA1A S2_31_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FA1A S2_31_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA1A S2_31_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA1A S2_31_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA1A S2_31_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA1A S2_31_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA1A S2_31_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA1A S2_31_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA1A S3_31_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\ab[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA1A S2_31_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), 
        .CO(\CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA1A S2_31_7 ( .A(\ab[31][7] ), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), 
        .CO(\CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA1A S2_31_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), 
        .CO(\CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA1A S2_31_4 ( .A(\ab[31][4] ), .B(\CARRYB[30][4] ), .CI(\SUMB[30][5] ), 
        .CO(\CARRYB[31][4] ), .S(\SUMB[31][4] ) );
  FA1A S2_31_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), 
        .CO(\CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA1A S2_31_3 ( .A(\ab[31][3] ), .B(\CARRYB[30][3] ), .CI(\SUMB[30][4] ), 
        .CO(\CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_30_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), 
        .CO(\CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA1A S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA1A S2_30_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), 
        .CO(\CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA1A S2_30_11 ( .A(\ab[30][11] ), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), 
        .CO(\CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA1A S2_30_12 ( .A(\ab[30][12] ), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), 
        .CO(\CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA1A S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), 
        .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA1A S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA1A S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA1A S2_30_16 ( .A(\ab[30][16] ), .B(\CARRYB[29][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA1A S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA1A S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA1A S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA1A S3_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\ab[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA1A S2_30_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), 
        .CO(\CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA1A S2_30_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), 
        .CO(\CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA1A S2_30_5 ( .A(\ab[30][5] ), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA1A S2_30_4 ( .A(\ab[30][4] ), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), 
        .CO(\CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA1A S2_30_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), 
        .CO(\CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA1A S2_30_3 ( .A(\ab[30][3] ), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), 
        .CO(\CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1A S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA1A S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA1A S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA1A S2_29_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA1A S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA1A S2_29_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA1A S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA1A S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA1A S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA1A S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA1A S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA1A S3_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\ab[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA1A S2_29_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1A S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA1A S2_29_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA1A S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1A S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1A S2_29_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA1A S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1A S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1A S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA1A S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA1A S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA1A S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA1A S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA1A S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA1A S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA1A S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA1A S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA1A S3_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\ab[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA1A S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1A S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1A S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1A S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1A S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1A S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1A S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1A S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA1A S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA1A S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA1A S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA1A S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA1A S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA1A S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA1A S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA1A S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA1A S3_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\ab[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA1A S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1A S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1A S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1A S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA1A S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1A S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA1A S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA1A S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1A S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA1A S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA1A S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA1A S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA1A S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA1A S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA1A S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA1A S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA1A S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA1A S3_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\ab[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA1A S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA1A S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA1A S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1A S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1A S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1A S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1A S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1A S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA1A S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA1A S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA1A S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA1A S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA1A S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA1A S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA1A S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA1A S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA1A S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA1A S3_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\ab[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA1A S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA1A S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA1A S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1A S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1A S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1A S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA1A S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1A S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA1A S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA1A S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA1A S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA1A S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA1A S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA1A S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA1A S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA1A S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA1A S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA1A S3_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\ab[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA1A S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1A S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1A S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA1A S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1A S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1A S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA1A S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA1A S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1A S2_23_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA1A S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA1A S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA1A S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA1A S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA1A S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA1A S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA1A S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA1A S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA1A S3_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\ab[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA1A S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1A S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1A S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1A S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1A S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1A S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1A S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA1A S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA1A S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA1A S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA1A S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA1A S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA1A S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA1A S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA1A S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA1A S3_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\ab[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA1A S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1A S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA1A S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA1A S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1A S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1A S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA1A S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA1A S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA1A S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA1A S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA1A S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA1A S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA1A S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA1A S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA1A S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA1A S3_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\ab[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA1A S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA1A S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA1A S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA1A S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA1A S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA1A S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA1A S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA1A S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA1A S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA1A S3_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\ab[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA1A S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA1A S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA1A S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA1A S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA1A S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA1A S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA1A S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA1A S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA1A S3_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\ab[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA1A S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA1A S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA1A S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA1A S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA1A S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA1A S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA1A S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA1A S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA1A S3_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\ab[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA1A S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA1A S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA1A S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA1A S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA1A S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA1A S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA1A S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA1A S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA1A S3_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\ab[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA1A S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA1A S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA1A S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA1A S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA1A S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA1A S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA1A S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA1A S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA1A S3_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\ab[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA1A S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA1A S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA1A S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA1A S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA1A S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA1A S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA1A S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA1A S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA1A S3_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\ab[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA1A S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA1A S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA1A S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA1A S3_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\ab[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA1A S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA1A S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA1A S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA1A S3_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\ab[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA1A S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA1A S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA1A S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA1A S3_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\ab[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA1A S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA1A S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA1A S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA1A S3_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\ab[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA1A S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA1A S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA1A S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA1A S3_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\ab[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA1A S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA1A S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA1A S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA1A S3_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\ab[8][21] ), .CO(
        \CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA1A S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA1A S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA1A S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA1A S3_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\ab[7][21] ), .CO(
        \CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA1A S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA1A S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA1A S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA1A S3_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\ab[6][21] ), .CO(
        \CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA1A S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA1A S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA1A S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA1A S3_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\ab[5][21] ), .CO(
        \CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA1A S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA1A S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA1A S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA1A S3_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\ab[4][21] ), .CO(
        \CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA1A S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA1A S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA1A S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA1A S3_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\ab[3][21] ), .CO(
        \CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA1A S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA1A S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA1A S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA1A S3_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\ab[2][21] ), .CO(
        \CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA1A S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA1A S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA1A S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA1A S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA1A S3_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\ab[1][21] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  EO U2 ( .A(\CARRYB[47][11] ), .B(\SUMB[47][12] ), .Z(\A1[57] ) );
  EO U3 ( .A(\CARRYB[47][10] ), .B(\SUMB[47][11] ), .Z(\A1[56] ) );
  EO U4 ( .A(\CARRYB[47][4] ), .B(\SUMB[47][5] ), .Z(\A1[50] ) );
  EO U5 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A1[48] ) );
  EO U6 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A1[51] ) );
  EO U7 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A1[54] ) );
  EO U8 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A1[52] ) );
  EO U9 ( .A(\CARRYB[47][7] ), .B(\SUMB[47][8] ), .Z(\A1[53] ) );
  EO U10 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A1[55] ) );
  EO U11 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A1[58] ) );
  EO U12 ( .A(\CARRYB[47][13] ), .B(\SUMB[47][14] ), .Z(\A1[59] ) );
  EO U13 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A1[60] ) );
  EO U14 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A1[47] ) );
  EO U15 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A1[49] ) );
  EO U16 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A1[61] ) );
  EO U17 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A1[62] ) );
  EO U18 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A1[64] ) );
  EO U19 ( .A(\CARRYB[47][17] ), .B(\SUMB[47][18] ), .Z(\A1[63] ) );
  EO U20 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A1[65] ) );
  EO U21 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A1[46] ) );
  EO U22 ( .A(\CARRYB[47][20] ), .B(\ab[47][21] ), .Z(\A1[66] ) );
  IVP U23 ( .A(B[20]), .Z(n6) );
  IVP U24 ( .A(B[19]), .Z(n7) );
  IVP U25 ( .A(B[18]), .Z(n8) );
  IVP U26 ( .A(B[17]), .Z(n9) );
  IVP U27 ( .A(B[21]), .Z(n5) );
  IVP U28 ( .A(B[0]), .Z(n13) );
  EO U29 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U30 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U31 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U32 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U33 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U34 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U35 ( .A(\ab[0][21] ), .B(\ab[1][20] ), .Z(\SUMB[1][20] ) );
  EO U36 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(\SUMB[1][19] ) );
  EO U37 ( .A(\ab[0][19] ), .B(\ab[1][18] ), .Z(\SUMB[1][18] ) );
  EO U38 ( .A(\ab[0][18] ), .B(\ab[1][17] ), .Z(\SUMB[1][17] ) );
  EO U39 ( .A(\ab[0][17] ), .B(\ab[1][16] ), .Z(\SUMB[1][16] ) );
  EO U40 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U41 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U42 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U43 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U44 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U45 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U46 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U47 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  IVP U48 ( .A(B[3]), .Z(n16) );
  IVP U49 ( .A(B[2]), .Z(n15) );
  IVP U50 ( .A(B[4]), .Z(n17) );
  IVP U51 ( .A(B[5]), .Z(n18) );
  IVP U52 ( .A(B[7]), .Z(n20) );
  IVP U53 ( .A(B[6]), .Z(n19) );
  IVP U54 ( .A(B[16]), .Z(n10) );
  IVP U55 ( .A(B[15]), .Z(n11) );
  IVP U56 ( .A(B[14]), .Z(n4) );
  IVP U57 ( .A(B[13]), .Z(n12) );
  IVP U58 ( .A(B[12]), .Z(n25) );
  IVP U59 ( .A(B[11]), .Z(n24) );
  IVP U60 ( .A(B[10]), .Z(n23) );
  IVP U61 ( .A(B[9]), .Z(n22) );
  IVP U62 ( .A(B[8]), .Z(n21) );
  IVP U63 ( .A(B[1]), .Z(n14) );
  IVP U64 ( .A(A[3]), .Z(n69) );
  IVP U65 ( .A(A[4]), .Z(n68) );
  IVP U66 ( .A(A[6]), .Z(n66) );
  IVP U67 ( .A(A[7]), .Z(n65) );
  IVP U68 ( .A(A[9]), .Z(n63) );
  IVP U69 ( .A(A[10]), .Z(n62) );
  IVP U70 ( .A(A[12]), .Z(n60) );
  IVP U71 ( .A(A[13]), .Z(n59) );
  IVP U72 ( .A(A[15]), .Z(n57) );
  IVP U73 ( .A(A[16]), .Z(n56) );
  IVP U74 ( .A(A[18]), .Z(n54) );
  IVP U75 ( .A(A[19]), .Z(n53) );
  IVP U76 ( .A(A[21]), .Z(n51) );
  IVP U77 ( .A(A[22]), .Z(n50) );
  IVP U78 ( .A(A[2]), .Z(n70) );
  IVP U79 ( .A(A[24]), .Z(n48) );
  IVP U80 ( .A(A[25]), .Z(n47) );
  IVP U81 ( .A(A[5]), .Z(n67) );
  IVP U82 ( .A(A[27]), .Z(n45) );
  IVP U83 ( .A(A[28]), .Z(n44) );
  IVP U84 ( .A(A[8]), .Z(n64) );
  IVP U85 ( .A(A[30]), .Z(n42) );
  IVP U86 ( .A(A[31]), .Z(n41) );
  IVP U87 ( .A(A[11]), .Z(n61) );
  IVP U88 ( .A(A[33]), .Z(n39) );
  IVP U89 ( .A(A[34]), .Z(n38) );
  IVP U90 ( .A(A[14]), .Z(n58) );
  IVP U91 ( .A(A[36]), .Z(n36) );
  IVP U92 ( .A(A[37]), .Z(n35) );
  IVP U93 ( .A(A[17]), .Z(n55) );
  IVP U94 ( .A(A[39]), .Z(n33) );
  IVP U95 ( .A(A[40]), .Z(n32) );
  IVP U96 ( .A(A[41]), .Z(n31) );
  IVP U97 ( .A(A[20]), .Z(n52) );
  IVP U98 ( .A(A[42]), .Z(n30) );
  IVP U99 ( .A(A[43]), .Z(n29) );
  IVP U100 ( .A(A[44]), .Z(n28) );
  IVP U101 ( .A(A[23]), .Z(n49) );
  IVP U102 ( .A(A[45]), .Z(n27) );
  IVP U103 ( .A(A[46]), .Z(n26) );
  IVP U104 ( .A(A[47]), .Z(n3) );
  IVP U105 ( .A(A[26]), .Z(n46) );
  IVP U106 ( .A(A[29]), .Z(n43) );
  IVP U107 ( .A(A[32]), .Z(n40) );
  IVP U108 ( .A(A[35]), .Z(n37) );
  IVP U109 ( .A(A[38]), .Z(n34) );
  IVP U110 ( .A(A[1]), .Z(n71) );
  IVP U111 ( .A(A[0]), .Z(n72) );
  EO U112 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  AN2P U113 ( .A(\CARRYB[47][0] ), .B(\SUMB[47][1] ), .Z(\A2[47] ) );
  AN2P U114 ( .A(\CARRYB[47][1] ), .B(\SUMB[47][2] ), .Z(\A2[48] ) );
  AN2P U115 ( .A(\CARRYB[47][2] ), .B(\SUMB[47][3] ), .Z(\A2[49] ) );
  AN2P U116 ( .A(\CARRYB[47][3] ), .B(\SUMB[47][4] ), .Z(\A2[50] ) );
  AN2P U117 ( .A(\CARRYB[47][4] ), .B(\SUMB[47][5] ), .Z(\A2[51] ) );
  AN2P U118 ( .A(\CARRYB[47][5] ), .B(\SUMB[47][6] ), .Z(\A2[52] ) );
  AN2P U119 ( .A(\CARRYB[47][6] ), .B(\SUMB[47][7] ), .Z(\A2[53] ) );
  AN2P U120 ( .A(\CARRYB[47][7] ), .B(\SUMB[47][8] ), .Z(\A2[54] ) );
  AN2P U121 ( .A(\CARRYB[47][8] ), .B(\SUMB[47][9] ), .Z(\A2[55] ) );
  AN2P U122 ( .A(\CARRYB[47][9] ), .B(\SUMB[47][10] ), .Z(\A2[56] ) );
  AN2P U123 ( .A(\CARRYB[47][10] ), .B(\SUMB[47][11] ), .Z(\A2[57] ) );
  AN2P U124 ( .A(\CARRYB[47][11] ), .B(\SUMB[47][12] ), .Z(\A2[58] ) );
  AN2P U125 ( .A(\CARRYB[47][12] ), .B(\SUMB[47][13] ), .Z(\A2[59] ) );
  AN2P U126 ( .A(\CARRYB[47][13] ), .B(\SUMB[47][14] ), .Z(\A2[60] ) );
  AN2P U127 ( .A(\CARRYB[47][14] ), .B(\SUMB[47][15] ), .Z(\A2[61] ) );
  AN2P U128 ( .A(\CARRYB[47][15] ), .B(\SUMB[47][16] ), .Z(\A2[62] ) );
  AN2P U129 ( .A(\CARRYB[47][16] ), .B(\SUMB[47][17] ), .Z(\A2[63] ) );
  AN2P U130 ( .A(\CARRYB[47][17] ), .B(\SUMB[47][18] ), .Z(\A2[64] ) );
  AN2P U131 ( .A(\CARRYB[47][18] ), .B(\SUMB[47][19] ), .Z(\A2[65] ) );
  AN2P U132 ( .A(\CARRYB[47][19] ), .B(\SUMB[47][20] ), .Z(\A2[66] ) );
  AN2P U133 ( .A(\CARRYB[47][20] ), .B(\ab[47][21] ), .Z(\A2[67] ) );
  AN2P U134 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U135 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U136 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U137 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U138 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U139 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U140 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U141 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U142 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U143 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U144 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U145 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U146 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U147 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U148 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U149 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\CARRYB[1][16] ) );
  AN2P U150 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\CARRYB[1][17] ) );
  AN2P U151 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\CARRYB[1][18] ) );
  AN2P U152 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\CARRYB[1][19] ) );
  AN2P U153 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\CARRYB[1][20] ) );
  NR2 U155 ( .A(n63), .B(n22), .Z(\ab[9][9] ) );
  NR2 U156 ( .A(n63), .B(n21), .Z(\ab[9][8] ) );
  NR2 U157 ( .A(n63), .B(n20), .Z(\ab[9][7] ) );
  NR2 U158 ( .A(n63), .B(n19), .Z(\ab[9][6] ) );
  NR2 U159 ( .A(n63), .B(n18), .Z(\ab[9][5] ) );
  NR2 U160 ( .A(n63), .B(n17), .Z(\ab[9][4] ) );
  NR2 U161 ( .A(n63), .B(n16), .Z(\ab[9][3] ) );
  NR2 U162 ( .A(n63), .B(n15), .Z(\ab[9][2] ) );
  NR2 U163 ( .A(n63), .B(n5), .Z(\ab[9][21] ) );
  NR2 U164 ( .A(n63), .B(n6), .Z(\ab[9][20] ) );
  NR2 U165 ( .A(n63), .B(n14), .Z(\ab[9][1] ) );
  NR2 U166 ( .A(n63), .B(n7), .Z(\ab[9][19] ) );
  NR2 U167 ( .A(n63), .B(n8), .Z(\ab[9][18] ) );
  NR2 U168 ( .A(n63), .B(n9), .Z(\ab[9][17] ) );
  NR2 U169 ( .A(n63), .B(n10), .Z(\ab[9][16] ) );
  NR2 U170 ( .A(n63), .B(n11), .Z(\ab[9][15] ) );
  NR2 U171 ( .A(n63), .B(n4), .Z(\ab[9][14] ) );
  NR2 U172 ( .A(n63), .B(n12), .Z(\ab[9][13] ) );
  NR2 U173 ( .A(n63), .B(n25), .Z(\ab[9][12] ) );
  NR2 U174 ( .A(n63), .B(n24), .Z(\ab[9][11] ) );
  NR2 U175 ( .A(n63), .B(n23), .Z(\ab[9][10] ) );
  NR2 U176 ( .A(n63), .B(n13), .Z(\ab[9][0] ) );
  NR2 U177 ( .A(n22), .B(n64), .Z(\ab[8][9] ) );
  NR2 U178 ( .A(n21), .B(n64), .Z(\ab[8][8] ) );
  NR2 U179 ( .A(n20), .B(n64), .Z(\ab[8][7] ) );
  NR2 U180 ( .A(n19), .B(n64), .Z(\ab[8][6] ) );
  NR2 U181 ( .A(n18), .B(n64), .Z(\ab[8][5] ) );
  NR2 U182 ( .A(n17), .B(n64), .Z(\ab[8][4] ) );
  NR2 U183 ( .A(n16), .B(n64), .Z(\ab[8][3] ) );
  NR2 U184 ( .A(n15), .B(n64), .Z(\ab[8][2] ) );
  NR2 U185 ( .A(n5), .B(n64), .Z(\ab[8][21] ) );
  NR2 U186 ( .A(n6), .B(n64), .Z(\ab[8][20] ) );
  NR2 U187 ( .A(n14), .B(n64), .Z(\ab[8][1] ) );
  NR2 U188 ( .A(n7), .B(n64), .Z(\ab[8][19] ) );
  NR2 U189 ( .A(n8), .B(n64), .Z(\ab[8][18] ) );
  NR2 U190 ( .A(n9), .B(n64), .Z(\ab[8][17] ) );
  NR2 U191 ( .A(n10), .B(n64), .Z(\ab[8][16] ) );
  NR2 U192 ( .A(n11), .B(n64), .Z(\ab[8][15] ) );
  NR2 U193 ( .A(n4), .B(n64), .Z(\ab[8][14] ) );
  NR2 U194 ( .A(n12), .B(n64), .Z(\ab[8][13] ) );
  NR2 U195 ( .A(n25), .B(n64), .Z(\ab[8][12] ) );
  NR2 U196 ( .A(n24), .B(n64), .Z(\ab[8][11] ) );
  NR2 U197 ( .A(n23), .B(n64), .Z(\ab[8][10] ) );
  NR2 U198 ( .A(n13), .B(n64), .Z(\ab[8][0] ) );
  NR2 U199 ( .A(n22), .B(n65), .Z(\ab[7][9] ) );
  NR2 U200 ( .A(n21), .B(n65), .Z(\ab[7][8] ) );
  NR2 U201 ( .A(n20), .B(n65), .Z(\ab[7][7] ) );
  NR2 U202 ( .A(n19), .B(n65), .Z(\ab[7][6] ) );
  NR2 U203 ( .A(n18), .B(n65), .Z(\ab[7][5] ) );
  NR2 U204 ( .A(n17), .B(n65), .Z(\ab[7][4] ) );
  NR2 U205 ( .A(n16), .B(n65), .Z(\ab[7][3] ) );
  NR2 U206 ( .A(n15), .B(n65), .Z(\ab[7][2] ) );
  NR2 U207 ( .A(n5), .B(n65), .Z(\ab[7][21] ) );
  NR2 U208 ( .A(n6), .B(n65), .Z(\ab[7][20] ) );
  NR2 U209 ( .A(n14), .B(n65), .Z(\ab[7][1] ) );
  NR2 U210 ( .A(n7), .B(n65), .Z(\ab[7][19] ) );
  NR2 U211 ( .A(n8), .B(n65), .Z(\ab[7][18] ) );
  NR2 U212 ( .A(n9), .B(n65), .Z(\ab[7][17] ) );
  NR2 U213 ( .A(n10), .B(n65), .Z(\ab[7][16] ) );
  NR2 U214 ( .A(n11), .B(n65), .Z(\ab[7][15] ) );
  NR2 U215 ( .A(n4), .B(n65), .Z(\ab[7][14] ) );
  NR2 U216 ( .A(n12), .B(n65), .Z(\ab[7][13] ) );
  NR2 U217 ( .A(n25), .B(n65), .Z(\ab[7][12] ) );
  NR2 U218 ( .A(n24), .B(n65), .Z(\ab[7][11] ) );
  NR2 U219 ( .A(n23), .B(n65), .Z(\ab[7][10] ) );
  NR2 U220 ( .A(n13), .B(n65), .Z(\ab[7][0] ) );
  NR2 U221 ( .A(n22), .B(n66), .Z(\ab[6][9] ) );
  NR2 U222 ( .A(n21), .B(n66), .Z(\ab[6][8] ) );
  NR2 U223 ( .A(n20), .B(n66), .Z(\ab[6][7] ) );
  NR2 U224 ( .A(n19), .B(n66), .Z(\ab[6][6] ) );
  NR2 U225 ( .A(n18), .B(n66), .Z(\ab[6][5] ) );
  NR2 U226 ( .A(n17), .B(n66), .Z(\ab[6][4] ) );
  NR2 U227 ( .A(n16), .B(n66), .Z(\ab[6][3] ) );
  NR2 U228 ( .A(n15), .B(n66), .Z(\ab[6][2] ) );
  NR2 U229 ( .A(n5), .B(n66), .Z(\ab[6][21] ) );
  NR2 U230 ( .A(n6), .B(n66), .Z(\ab[6][20] ) );
  NR2 U231 ( .A(n14), .B(n66), .Z(\ab[6][1] ) );
  NR2 U232 ( .A(n7), .B(n66), .Z(\ab[6][19] ) );
  NR2 U233 ( .A(n8), .B(n66), .Z(\ab[6][18] ) );
  NR2 U234 ( .A(n9), .B(n66), .Z(\ab[6][17] ) );
  NR2 U235 ( .A(n10), .B(n66), .Z(\ab[6][16] ) );
  NR2 U236 ( .A(n11), .B(n66), .Z(\ab[6][15] ) );
  NR2 U237 ( .A(n4), .B(n66), .Z(\ab[6][14] ) );
  NR2 U238 ( .A(n12), .B(n66), .Z(\ab[6][13] ) );
  NR2 U239 ( .A(n25), .B(n66), .Z(\ab[6][12] ) );
  NR2 U240 ( .A(n24), .B(n66), .Z(\ab[6][11] ) );
  NR2 U241 ( .A(n23), .B(n66), .Z(\ab[6][10] ) );
  NR2 U242 ( .A(n13), .B(n66), .Z(\ab[6][0] ) );
  NR2 U243 ( .A(n22), .B(n67), .Z(\ab[5][9] ) );
  NR2 U244 ( .A(n21), .B(n67), .Z(\ab[5][8] ) );
  NR2 U245 ( .A(n20), .B(n67), .Z(\ab[5][7] ) );
  NR2 U246 ( .A(n19), .B(n67), .Z(\ab[5][6] ) );
  NR2 U247 ( .A(n18), .B(n67), .Z(\ab[5][5] ) );
  NR2 U248 ( .A(n17), .B(n67), .Z(\ab[5][4] ) );
  NR2 U249 ( .A(n16), .B(n67), .Z(\ab[5][3] ) );
  NR2 U250 ( .A(n15), .B(n67), .Z(\ab[5][2] ) );
  NR2 U251 ( .A(n5), .B(n67), .Z(\ab[5][21] ) );
  NR2 U252 ( .A(n6), .B(n67), .Z(\ab[5][20] ) );
  NR2 U253 ( .A(n14), .B(n67), .Z(\ab[5][1] ) );
  NR2 U254 ( .A(n7), .B(n67), .Z(\ab[5][19] ) );
  NR2 U255 ( .A(n8), .B(n67), .Z(\ab[5][18] ) );
  NR2 U256 ( .A(n9), .B(n67), .Z(\ab[5][17] ) );
  NR2 U257 ( .A(n10), .B(n67), .Z(\ab[5][16] ) );
  NR2 U258 ( .A(n11), .B(n67), .Z(\ab[5][15] ) );
  NR2 U259 ( .A(n4), .B(n67), .Z(\ab[5][14] ) );
  NR2 U260 ( .A(n12), .B(n67), .Z(\ab[5][13] ) );
  NR2 U261 ( .A(n25), .B(n67), .Z(\ab[5][12] ) );
  NR2 U262 ( .A(n24), .B(n67), .Z(\ab[5][11] ) );
  NR2 U263 ( .A(n23), .B(n67), .Z(\ab[5][10] ) );
  NR2 U264 ( .A(n13), .B(n67), .Z(\ab[5][0] ) );
  NR2 U265 ( .A(n22), .B(n68), .Z(\ab[4][9] ) );
  NR2 U266 ( .A(n21), .B(n68), .Z(\ab[4][8] ) );
  NR2 U267 ( .A(n20), .B(n68), .Z(\ab[4][7] ) );
  NR2 U268 ( .A(n19), .B(n68), .Z(\ab[4][6] ) );
  NR2 U269 ( .A(n18), .B(n68), .Z(\ab[4][5] ) );
  NR2 U270 ( .A(n17), .B(n68), .Z(\ab[4][4] ) );
  NR2 U271 ( .A(n16), .B(n68), .Z(\ab[4][3] ) );
  NR2 U272 ( .A(n15), .B(n68), .Z(\ab[4][2] ) );
  NR2 U273 ( .A(n5), .B(n68), .Z(\ab[4][21] ) );
  NR2 U274 ( .A(n6), .B(n68), .Z(\ab[4][20] ) );
  NR2 U275 ( .A(n14), .B(n68), .Z(\ab[4][1] ) );
  NR2 U276 ( .A(n7), .B(n68), .Z(\ab[4][19] ) );
  NR2 U277 ( .A(n8), .B(n68), .Z(\ab[4][18] ) );
  NR2 U278 ( .A(n9), .B(n68), .Z(\ab[4][17] ) );
  NR2 U279 ( .A(n10), .B(n68), .Z(\ab[4][16] ) );
  NR2 U280 ( .A(n11), .B(n68), .Z(\ab[4][15] ) );
  NR2 U281 ( .A(n4), .B(n68), .Z(\ab[4][14] ) );
  NR2 U282 ( .A(n12), .B(n68), .Z(\ab[4][13] ) );
  NR2 U283 ( .A(n25), .B(n68), .Z(\ab[4][12] ) );
  NR2 U284 ( .A(n24), .B(n68), .Z(\ab[4][11] ) );
  NR2 U285 ( .A(n23), .B(n68), .Z(\ab[4][10] ) );
  NR2 U286 ( .A(n13), .B(n68), .Z(\ab[4][0] ) );
  NR2 U287 ( .A(n22), .B(n3), .Z(\ab[47][9] ) );
  NR2 U288 ( .A(n21), .B(n3), .Z(\ab[47][8] ) );
  NR2 U289 ( .A(n20), .B(n3), .Z(\ab[47][7] ) );
  NR2 U290 ( .A(n19), .B(n3), .Z(\ab[47][6] ) );
  NR2 U291 ( .A(n18), .B(n3), .Z(\ab[47][5] ) );
  NR2 U292 ( .A(n17), .B(n3), .Z(\ab[47][4] ) );
  NR2 U293 ( .A(n16), .B(n3), .Z(\ab[47][3] ) );
  NR2 U294 ( .A(n15), .B(n3), .Z(\ab[47][2] ) );
  NR2 U295 ( .A(n5), .B(n3), .Z(\ab[47][21] ) );
  NR2 U296 ( .A(n6), .B(n3), .Z(\ab[47][20] ) );
  NR2 U297 ( .A(n14), .B(n3), .Z(\ab[47][1] ) );
  NR2 U298 ( .A(n7), .B(n3), .Z(\ab[47][19] ) );
  NR2 U299 ( .A(n8), .B(n3), .Z(\ab[47][18] ) );
  NR2 U300 ( .A(n9), .B(n3), .Z(\ab[47][17] ) );
  NR2 U301 ( .A(n10), .B(n3), .Z(\ab[47][16] ) );
  NR2 U302 ( .A(n11), .B(n3), .Z(\ab[47][15] ) );
  NR2 U303 ( .A(n4), .B(n3), .Z(\ab[47][14] ) );
  NR2 U304 ( .A(n12), .B(n3), .Z(\ab[47][13] ) );
  NR2 U305 ( .A(n25), .B(n3), .Z(\ab[47][12] ) );
  NR2 U306 ( .A(n24), .B(n3), .Z(\ab[47][11] ) );
  NR2 U307 ( .A(n23), .B(n3), .Z(\ab[47][10] ) );
  NR2 U308 ( .A(n13), .B(n3), .Z(\ab[47][0] ) );
  NR2 U309 ( .A(n22), .B(n26), .Z(\ab[46][9] ) );
  NR2 U310 ( .A(n21), .B(n26), .Z(\ab[46][8] ) );
  NR2 U311 ( .A(n20), .B(n26), .Z(\ab[46][7] ) );
  NR2 U312 ( .A(n19), .B(n26), .Z(\ab[46][6] ) );
  NR2 U313 ( .A(n18), .B(n26), .Z(\ab[46][5] ) );
  NR2 U314 ( .A(n17), .B(n26), .Z(\ab[46][4] ) );
  NR2 U315 ( .A(n16), .B(n26), .Z(\ab[46][3] ) );
  NR2 U316 ( .A(n15), .B(n26), .Z(\ab[46][2] ) );
  NR2 U317 ( .A(n5), .B(n26), .Z(\ab[46][21] ) );
  NR2 U318 ( .A(n6), .B(n26), .Z(\ab[46][20] ) );
  NR2 U319 ( .A(n14), .B(n26), .Z(\ab[46][1] ) );
  NR2 U320 ( .A(n7), .B(n26), .Z(\ab[46][19] ) );
  NR2 U321 ( .A(n8), .B(n26), .Z(\ab[46][18] ) );
  NR2 U322 ( .A(n9), .B(n26), .Z(\ab[46][17] ) );
  NR2 U323 ( .A(n10), .B(n26), .Z(\ab[46][16] ) );
  NR2 U324 ( .A(n11), .B(n26), .Z(\ab[46][15] ) );
  NR2 U325 ( .A(n4), .B(n26), .Z(\ab[46][14] ) );
  NR2 U326 ( .A(n12), .B(n26), .Z(\ab[46][13] ) );
  NR2 U327 ( .A(n25), .B(n26), .Z(\ab[46][12] ) );
  NR2 U328 ( .A(n24), .B(n26), .Z(\ab[46][11] ) );
  NR2 U329 ( .A(n23), .B(n26), .Z(\ab[46][10] ) );
  NR2 U330 ( .A(n13), .B(n26), .Z(\ab[46][0] ) );
  NR2 U331 ( .A(n22), .B(n27), .Z(\ab[45][9] ) );
  NR2 U332 ( .A(n21), .B(n27), .Z(\ab[45][8] ) );
  NR2 U333 ( .A(n20), .B(n27), .Z(\ab[45][7] ) );
  NR2 U334 ( .A(n19), .B(n27), .Z(\ab[45][6] ) );
  NR2 U335 ( .A(n18), .B(n27), .Z(\ab[45][5] ) );
  NR2 U336 ( .A(n17), .B(n27), .Z(\ab[45][4] ) );
  NR2 U337 ( .A(n16), .B(n27), .Z(\ab[45][3] ) );
  NR2 U338 ( .A(n15), .B(n27), .Z(\ab[45][2] ) );
  NR2 U339 ( .A(n5), .B(n27), .Z(\ab[45][21] ) );
  NR2 U340 ( .A(n6), .B(n27), .Z(\ab[45][20] ) );
  NR2 U341 ( .A(n14), .B(n27), .Z(\ab[45][1] ) );
  NR2 U342 ( .A(n7), .B(n27), .Z(\ab[45][19] ) );
  NR2 U343 ( .A(n8), .B(n27), .Z(\ab[45][18] ) );
  NR2 U344 ( .A(n9), .B(n27), .Z(\ab[45][17] ) );
  NR2 U345 ( .A(n10), .B(n27), .Z(\ab[45][16] ) );
  NR2 U346 ( .A(n11), .B(n27), .Z(\ab[45][15] ) );
  NR2 U347 ( .A(n4), .B(n27), .Z(\ab[45][14] ) );
  NR2 U348 ( .A(n12), .B(n27), .Z(\ab[45][13] ) );
  NR2 U349 ( .A(n25), .B(n27), .Z(\ab[45][12] ) );
  NR2 U350 ( .A(n24), .B(n27), .Z(\ab[45][11] ) );
  NR2 U351 ( .A(n23), .B(n27), .Z(\ab[45][10] ) );
  NR2 U352 ( .A(n13), .B(n27), .Z(\ab[45][0] ) );
  NR2 U353 ( .A(n22), .B(n28), .Z(\ab[44][9] ) );
  NR2 U354 ( .A(n21), .B(n28), .Z(\ab[44][8] ) );
  NR2 U355 ( .A(n20), .B(n28), .Z(\ab[44][7] ) );
  NR2 U356 ( .A(n19), .B(n28), .Z(\ab[44][6] ) );
  NR2 U357 ( .A(n18), .B(n28), .Z(\ab[44][5] ) );
  NR2 U358 ( .A(n17), .B(n28), .Z(\ab[44][4] ) );
  NR2 U359 ( .A(n16), .B(n28), .Z(\ab[44][3] ) );
  NR2 U360 ( .A(n15), .B(n28), .Z(\ab[44][2] ) );
  NR2 U361 ( .A(n5), .B(n28), .Z(\ab[44][21] ) );
  NR2 U362 ( .A(n6), .B(n28), .Z(\ab[44][20] ) );
  NR2 U363 ( .A(n14), .B(n28), .Z(\ab[44][1] ) );
  NR2 U364 ( .A(n7), .B(n28), .Z(\ab[44][19] ) );
  NR2 U365 ( .A(n8), .B(n28), .Z(\ab[44][18] ) );
  NR2 U366 ( .A(n9), .B(n28), .Z(\ab[44][17] ) );
  NR2 U367 ( .A(n10), .B(n28), .Z(\ab[44][16] ) );
  NR2 U368 ( .A(n11), .B(n28), .Z(\ab[44][15] ) );
  NR2 U369 ( .A(n4), .B(n28), .Z(\ab[44][14] ) );
  NR2 U370 ( .A(n12), .B(n28), .Z(\ab[44][13] ) );
  NR2 U371 ( .A(n25), .B(n28), .Z(\ab[44][12] ) );
  NR2 U372 ( .A(n24), .B(n28), .Z(\ab[44][11] ) );
  NR2 U373 ( .A(n23), .B(n28), .Z(\ab[44][10] ) );
  NR2 U374 ( .A(n13), .B(n28), .Z(\ab[44][0] ) );
  NR2 U375 ( .A(n22), .B(n29), .Z(\ab[43][9] ) );
  NR2 U376 ( .A(n21), .B(n29), .Z(\ab[43][8] ) );
  NR2 U377 ( .A(n20), .B(n29), .Z(\ab[43][7] ) );
  NR2 U378 ( .A(n19), .B(n29), .Z(\ab[43][6] ) );
  NR2 U379 ( .A(n18), .B(n29), .Z(\ab[43][5] ) );
  NR2 U380 ( .A(n17), .B(n29), .Z(\ab[43][4] ) );
  NR2 U381 ( .A(n16), .B(n29), .Z(\ab[43][3] ) );
  NR2 U382 ( .A(n15), .B(n29), .Z(\ab[43][2] ) );
  NR2 U383 ( .A(n5), .B(n29), .Z(\ab[43][21] ) );
  NR2 U384 ( .A(n6), .B(n29), .Z(\ab[43][20] ) );
  NR2 U385 ( .A(n14), .B(n29), .Z(\ab[43][1] ) );
  NR2 U386 ( .A(n7), .B(n29), .Z(\ab[43][19] ) );
  NR2 U387 ( .A(n8), .B(n29), .Z(\ab[43][18] ) );
  NR2 U388 ( .A(n9), .B(n29), .Z(\ab[43][17] ) );
  NR2 U389 ( .A(n10), .B(n29), .Z(\ab[43][16] ) );
  NR2 U390 ( .A(n11), .B(n29), .Z(\ab[43][15] ) );
  NR2 U391 ( .A(n4), .B(n29), .Z(\ab[43][14] ) );
  NR2 U392 ( .A(n12), .B(n29), .Z(\ab[43][13] ) );
  NR2 U393 ( .A(n25), .B(n29), .Z(\ab[43][12] ) );
  NR2 U394 ( .A(n24), .B(n29), .Z(\ab[43][11] ) );
  NR2 U395 ( .A(n23), .B(n29), .Z(\ab[43][10] ) );
  NR2 U396 ( .A(n13), .B(n29), .Z(\ab[43][0] ) );
  NR2 U397 ( .A(n22), .B(n30), .Z(\ab[42][9] ) );
  NR2 U398 ( .A(n21), .B(n30), .Z(\ab[42][8] ) );
  NR2 U399 ( .A(n20), .B(n30), .Z(\ab[42][7] ) );
  NR2 U400 ( .A(n19), .B(n30), .Z(\ab[42][6] ) );
  NR2 U401 ( .A(n18), .B(n30), .Z(\ab[42][5] ) );
  NR2 U402 ( .A(n17), .B(n30), .Z(\ab[42][4] ) );
  NR2 U403 ( .A(n16), .B(n30), .Z(\ab[42][3] ) );
  NR2 U404 ( .A(n15), .B(n30), .Z(\ab[42][2] ) );
  NR2 U405 ( .A(n5), .B(n30), .Z(\ab[42][21] ) );
  NR2 U406 ( .A(n6), .B(n30), .Z(\ab[42][20] ) );
  NR2 U407 ( .A(n14), .B(n30), .Z(\ab[42][1] ) );
  NR2 U408 ( .A(n7), .B(n30), .Z(\ab[42][19] ) );
  NR2 U409 ( .A(n8), .B(n30), .Z(\ab[42][18] ) );
  NR2 U410 ( .A(n9), .B(n30), .Z(\ab[42][17] ) );
  NR2 U411 ( .A(n10), .B(n30), .Z(\ab[42][16] ) );
  NR2 U412 ( .A(n11), .B(n30), .Z(\ab[42][15] ) );
  NR2 U413 ( .A(n4), .B(n30), .Z(\ab[42][14] ) );
  NR2 U414 ( .A(n12), .B(n30), .Z(\ab[42][13] ) );
  NR2 U415 ( .A(n25), .B(n30), .Z(\ab[42][12] ) );
  NR2 U416 ( .A(n24), .B(n30), .Z(\ab[42][11] ) );
  NR2 U417 ( .A(n23), .B(n30), .Z(\ab[42][10] ) );
  NR2 U418 ( .A(n13), .B(n30), .Z(\ab[42][0] ) );
  NR2 U419 ( .A(n22), .B(n31), .Z(\ab[41][9] ) );
  NR2 U420 ( .A(n21), .B(n31), .Z(\ab[41][8] ) );
  NR2 U421 ( .A(n20), .B(n31), .Z(\ab[41][7] ) );
  NR2 U422 ( .A(n19), .B(n31), .Z(\ab[41][6] ) );
  NR2 U423 ( .A(n18), .B(n31), .Z(\ab[41][5] ) );
  NR2 U424 ( .A(n17), .B(n31), .Z(\ab[41][4] ) );
  NR2 U425 ( .A(n16), .B(n31), .Z(\ab[41][3] ) );
  NR2 U426 ( .A(n15), .B(n31), .Z(\ab[41][2] ) );
  NR2 U427 ( .A(n5), .B(n31), .Z(\ab[41][21] ) );
  NR2 U428 ( .A(n6), .B(n31), .Z(\ab[41][20] ) );
  NR2 U429 ( .A(n14), .B(n31), .Z(\ab[41][1] ) );
  NR2 U430 ( .A(n7), .B(n31), .Z(\ab[41][19] ) );
  NR2 U431 ( .A(n8), .B(n31), .Z(\ab[41][18] ) );
  NR2 U432 ( .A(n9), .B(n31), .Z(\ab[41][17] ) );
  NR2 U433 ( .A(n10), .B(n31), .Z(\ab[41][16] ) );
  NR2 U434 ( .A(n11), .B(n31), .Z(\ab[41][15] ) );
  NR2 U435 ( .A(n4), .B(n31), .Z(\ab[41][14] ) );
  NR2 U436 ( .A(n12), .B(n31), .Z(\ab[41][13] ) );
  NR2 U437 ( .A(n25), .B(n31), .Z(\ab[41][12] ) );
  NR2 U438 ( .A(n24), .B(n31), .Z(\ab[41][11] ) );
  NR2 U439 ( .A(n23), .B(n31), .Z(\ab[41][10] ) );
  NR2 U440 ( .A(n13), .B(n31), .Z(\ab[41][0] ) );
  NR2 U441 ( .A(n22), .B(n32), .Z(\ab[40][9] ) );
  NR2 U442 ( .A(n21), .B(n32), .Z(\ab[40][8] ) );
  NR2 U443 ( .A(n20), .B(n32), .Z(\ab[40][7] ) );
  NR2 U444 ( .A(n19), .B(n32), .Z(\ab[40][6] ) );
  NR2 U445 ( .A(n18), .B(n32), .Z(\ab[40][5] ) );
  NR2 U446 ( .A(n17), .B(n32), .Z(\ab[40][4] ) );
  NR2 U447 ( .A(n16), .B(n32), .Z(\ab[40][3] ) );
  NR2 U448 ( .A(n15), .B(n32), .Z(\ab[40][2] ) );
  NR2 U449 ( .A(n5), .B(n32), .Z(\ab[40][21] ) );
  NR2 U450 ( .A(n6), .B(n32), .Z(\ab[40][20] ) );
  NR2 U451 ( .A(n14), .B(n32), .Z(\ab[40][1] ) );
  NR2 U452 ( .A(n7), .B(n32), .Z(\ab[40][19] ) );
  NR2 U453 ( .A(n8), .B(n32), .Z(\ab[40][18] ) );
  NR2 U454 ( .A(n9), .B(n32), .Z(\ab[40][17] ) );
  NR2 U455 ( .A(n10), .B(n32), .Z(\ab[40][16] ) );
  NR2 U456 ( .A(n11), .B(n32), .Z(\ab[40][15] ) );
  NR2 U457 ( .A(n4), .B(n32), .Z(\ab[40][14] ) );
  NR2 U458 ( .A(n12), .B(n32), .Z(\ab[40][13] ) );
  NR2 U459 ( .A(n25), .B(n32), .Z(\ab[40][12] ) );
  NR2 U460 ( .A(n24), .B(n32), .Z(\ab[40][11] ) );
  NR2 U461 ( .A(n23), .B(n32), .Z(\ab[40][10] ) );
  NR2 U462 ( .A(n13), .B(n32), .Z(\ab[40][0] ) );
  NR2 U463 ( .A(n22), .B(n69), .Z(\ab[3][9] ) );
  NR2 U464 ( .A(n21), .B(n69), .Z(\ab[3][8] ) );
  NR2 U465 ( .A(n20), .B(n69), .Z(\ab[3][7] ) );
  NR2 U466 ( .A(n19), .B(n69), .Z(\ab[3][6] ) );
  NR2 U467 ( .A(n18), .B(n69), .Z(\ab[3][5] ) );
  NR2 U468 ( .A(n17), .B(n69), .Z(\ab[3][4] ) );
  NR2 U469 ( .A(n16), .B(n69), .Z(\ab[3][3] ) );
  NR2 U470 ( .A(n15), .B(n69), .Z(\ab[3][2] ) );
  NR2 U471 ( .A(n5), .B(n69), .Z(\ab[3][21] ) );
  NR2 U472 ( .A(n6), .B(n69), .Z(\ab[3][20] ) );
  NR2 U473 ( .A(n14), .B(n69), .Z(\ab[3][1] ) );
  NR2 U474 ( .A(n7), .B(n69), .Z(\ab[3][19] ) );
  NR2 U475 ( .A(n8), .B(n69), .Z(\ab[3][18] ) );
  NR2 U476 ( .A(n9), .B(n69), .Z(\ab[3][17] ) );
  NR2 U477 ( .A(n10), .B(n69), .Z(\ab[3][16] ) );
  NR2 U478 ( .A(n11), .B(n69), .Z(\ab[3][15] ) );
  NR2 U479 ( .A(n4), .B(n69), .Z(\ab[3][14] ) );
  NR2 U480 ( .A(n12), .B(n69), .Z(\ab[3][13] ) );
  NR2 U481 ( .A(n25), .B(n69), .Z(\ab[3][12] ) );
  NR2 U482 ( .A(n24), .B(n69), .Z(\ab[3][11] ) );
  NR2 U483 ( .A(n23), .B(n69), .Z(\ab[3][10] ) );
  NR2 U484 ( .A(n13), .B(n69), .Z(\ab[3][0] ) );
  NR2 U485 ( .A(n22), .B(n33), .Z(\ab[39][9] ) );
  NR2 U486 ( .A(n21), .B(n33), .Z(\ab[39][8] ) );
  NR2 U487 ( .A(n20), .B(n33), .Z(\ab[39][7] ) );
  NR2 U488 ( .A(n19), .B(n33), .Z(\ab[39][6] ) );
  NR2 U489 ( .A(n18), .B(n33), .Z(\ab[39][5] ) );
  NR2 U490 ( .A(n17), .B(n33), .Z(\ab[39][4] ) );
  NR2 U491 ( .A(n16), .B(n33), .Z(\ab[39][3] ) );
  NR2 U492 ( .A(n15), .B(n33), .Z(\ab[39][2] ) );
  NR2 U493 ( .A(n5), .B(n33), .Z(\ab[39][21] ) );
  NR2 U494 ( .A(n6), .B(n33), .Z(\ab[39][20] ) );
  NR2 U495 ( .A(n14), .B(n33), .Z(\ab[39][1] ) );
  NR2 U496 ( .A(n7), .B(n33), .Z(\ab[39][19] ) );
  NR2 U497 ( .A(n8), .B(n33), .Z(\ab[39][18] ) );
  NR2 U498 ( .A(n9), .B(n33), .Z(\ab[39][17] ) );
  NR2 U499 ( .A(n10), .B(n33), .Z(\ab[39][16] ) );
  NR2 U500 ( .A(n11), .B(n33), .Z(\ab[39][15] ) );
  NR2 U501 ( .A(n4), .B(n33), .Z(\ab[39][14] ) );
  NR2 U502 ( .A(n12), .B(n33), .Z(\ab[39][13] ) );
  NR2 U503 ( .A(n25), .B(n33), .Z(\ab[39][12] ) );
  NR2 U504 ( .A(n24), .B(n33), .Z(\ab[39][11] ) );
  NR2 U505 ( .A(n23), .B(n33), .Z(\ab[39][10] ) );
  NR2 U506 ( .A(n13), .B(n33), .Z(\ab[39][0] ) );
  NR2 U507 ( .A(n22), .B(n34), .Z(\ab[38][9] ) );
  NR2 U508 ( .A(n21), .B(n34), .Z(\ab[38][8] ) );
  NR2 U509 ( .A(n20), .B(n34), .Z(\ab[38][7] ) );
  NR2 U510 ( .A(n19), .B(n34), .Z(\ab[38][6] ) );
  NR2 U511 ( .A(n18), .B(n34), .Z(\ab[38][5] ) );
  NR2 U512 ( .A(n17), .B(n34), .Z(\ab[38][4] ) );
  NR2 U513 ( .A(n16), .B(n34), .Z(\ab[38][3] ) );
  NR2 U514 ( .A(n15), .B(n34), .Z(\ab[38][2] ) );
  NR2 U515 ( .A(n5), .B(n34), .Z(\ab[38][21] ) );
  NR2 U516 ( .A(n6), .B(n34), .Z(\ab[38][20] ) );
  NR2 U517 ( .A(n14), .B(n34), .Z(\ab[38][1] ) );
  NR2 U518 ( .A(n7), .B(n34), .Z(\ab[38][19] ) );
  NR2 U519 ( .A(n8), .B(n34), .Z(\ab[38][18] ) );
  NR2 U520 ( .A(n9), .B(n34), .Z(\ab[38][17] ) );
  NR2 U521 ( .A(n10), .B(n34), .Z(\ab[38][16] ) );
  NR2 U522 ( .A(n11), .B(n34), .Z(\ab[38][15] ) );
  NR2 U523 ( .A(n4), .B(n34), .Z(\ab[38][14] ) );
  NR2 U524 ( .A(n12), .B(n34), .Z(\ab[38][13] ) );
  NR2 U525 ( .A(n25), .B(n34), .Z(\ab[38][12] ) );
  NR2 U526 ( .A(n24), .B(n34), .Z(\ab[38][11] ) );
  NR2 U527 ( .A(n23), .B(n34), .Z(\ab[38][10] ) );
  NR2 U528 ( .A(n13), .B(n34), .Z(\ab[38][0] ) );
  NR2 U529 ( .A(n22), .B(n35), .Z(\ab[37][9] ) );
  NR2 U530 ( .A(n21), .B(n35), .Z(\ab[37][8] ) );
  NR2 U531 ( .A(n20), .B(n35), .Z(\ab[37][7] ) );
  NR2 U532 ( .A(n19), .B(n35), .Z(\ab[37][6] ) );
  NR2 U533 ( .A(n18), .B(n35), .Z(\ab[37][5] ) );
  NR2 U534 ( .A(n17), .B(n35), .Z(\ab[37][4] ) );
  NR2 U535 ( .A(n16), .B(n35), .Z(\ab[37][3] ) );
  NR2 U536 ( .A(n15), .B(n35), .Z(\ab[37][2] ) );
  NR2 U537 ( .A(n5), .B(n35), .Z(\ab[37][21] ) );
  NR2 U538 ( .A(n6), .B(n35), .Z(\ab[37][20] ) );
  NR2 U539 ( .A(n14), .B(n35), .Z(\ab[37][1] ) );
  NR2 U540 ( .A(n7), .B(n35), .Z(\ab[37][19] ) );
  NR2 U541 ( .A(n8), .B(n35), .Z(\ab[37][18] ) );
  NR2 U542 ( .A(n9), .B(n35), .Z(\ab[37][17] ) );
  NR2 U543 ( .A(n10), .B(n35), .Z(\ab[37][16] ) );
  NR2 U544 ( .A(n11), .B(n35), .Z(\ab[37][15] ) );
  NR2 U545 ( .A(n4), .B(n35), .Z(\ab[37][14] ) );
  NR2 U546 ( .A(n12), .B(n35), .Z(\ab[37][13] ) );
  NR2 U547 ( .A(n25), .B(n35), .Z(\ab[37][12] ) );
  NR2 U548 ( .A(n24), .B(n35), .Z(\ab[37][11] ) );
  NR2 U549 ( .A(n23), .B(n35), .Z(\ab[37][10] ) );
  NR2 U550 ( .A(n13), .B(n35), .Z(\ab[37][0] ) );
  NR2 U551 ( .A(n22), .B(n36), .Z(\ab[36][9] ) );
  NR2 U552 ( .A(n21), .B(n36), .Z(\ab[36][8] ) );
  NR2 U553 ( .A(n20), .B(n36), .Z(\ab[36][7] ) );
  NR2 U554 ( .A(n19), .B(n36), .Z(\ab[36][6] ) );
  NR2 U555 ( .A(n18), .B(n36), .Z(\ab[36][5] ) );
  NR2 U556 ( .A(n17), .B(n36), .Z(\ab[36][4] ) );
  NR2 U557 ( .A(n16), .B(n36), .Z(\ab[36][3] ) );
  NR2 U558 ( .A(n15), .B(n36), .Z(\ab[36][2] ) );
  NR2 U559 ( .A(n5), .B(n36), .Z(\ab[36][21] ) );
  NR2 U560 ( .A(n6), .B(n36), .Z(\ab[36][20] ) );
  NR2 U561 ( .A(n14), .B(n36), .Z(\ab[36][1] ) );
  NR2 U562 ( .A(n7), .B(n36), .Z(\ab[36][19] ) );
  NR2 U563 ( .A(n8), .B(n36), .Z(\ab[36][18] ) );
  NR2 U564 ( .A(n9), .B(n36), .Z(\ab[36][17] ) );
  NR2 U565 ( .A(n10), .B(n36), .Z(\ab[36][16] ) );
  NR2 U566 ( .A(n11), .B(n36), .Z(\ab[36][15] ) );
  NR2 U567 ( .A(n4), .B(n36), .Z(\ab[36][14] ) );
  NR2 U568 ( .A(n12), .B(n36), .Z(\ab[36][13] ) );
  NR2 U569 ( .A(n25), .B(n36), .Z(\ab[36][12] ) );
  NR2 U570 ( .A(n24), .B(n36), .Z(\ab[36][11] ) );
  NR2 U571 ( .A(n23), .B(n36), .Z(\ab[36][10] ) );
  NR2 U572 ( .A(n13), .B(n36), .Z(\ab[36][0] ) );
  NR2 U573 ( .A(n22), .B(n37), .Z(\ab[35][9] ) );
  NR2 U574 ( .A(n21), .B(n37), .Z(\ab[35][8] ) );
  NR2 U575 ( .A(n20), .B(n37), .Z(\ab[35][7] ) );
  NR2 U576 ( .A(n19), .B(n37), .Z(\ab[35][6] ) );
  NR2 U577 ( .A(n18), .B(n37), .Z(\ab[35][5] ) );
  NR2 U578 ( .A(n17), .B(n37), .Z(\ab[35][4] ) );
  NR2 U579 ( .A(n16), .B(n37), .Z(\ab[35][3] ) );
  NR2 U580 ( .A(n15), .B(n37), .Z(\ab[35][2] ) );
  NR2 U581 ( .A(n5), .B(n37), .Z(\ab[35][21] ) );
  NR2 U582 ( .A(n6), .B(n37), .Z(\ab[35][20] ) );
  NR2 U583 ( .A(n14), .B(n37), .Z(\ab[35][1] ) );
  NR2 U584 ( .A(n7), .B(n37), .Z(\ab[35][19] ) );
  NR2 U585 ( .A(n8), .B(n37), .Z(\ab[35][18] ) );
  NR2 U586 ( .A(n9), .B(n37), .Z(\ab[35][17] ) );
  NR2 U587 ( .A(n10), .B(n37), .Z(\ab[35][16] ) );
  NR2 U588 ( .A(n11), .B(n37), .Z(\ab[35][15] ) );
  NR2 U589 ( .A(n4), .B(n37), .Z(\ab[35][14] ) );
  NR2 U590 ( .A(n12), .B(n37), .Z(\ab[35][13] ) );
  NR2 U591 ( .A(n25), .B(n37), .Z(\ab[35][12] ) );
  NR2 U592 ( .A(n24), .B(n37), .Z(\ab[35][11] ) );
  NR2 U593 ( .A(n23), .B(n37), .Z(\ab[35][10] ) );
  NR2 U594 ( .A(n13), .B(n37), .Z(\ab[35][0] ) );
  NR2 U595 ( .A(n22), .B(n38), .Z(\ab[34][9] ) );
  NR2 U596 ( .A(n21), .B(n38), .Z(\ab[34][8] ) );
  NR2 U597 ( .A(n20), .B(n38), .Z(\ab[34][7] ) );
  NR2 U598 ( .A(n19), .B(n38), .Z(\ab[34][6] ) );
  NR2 U599 ( .A(n18), .B(n38), .Z(\ab[34][5] ) );
  NR2 U600 ( .A(n17), .B(n38), .Z(\ab[34][4] ) );
  NR2 U601 ( .A(n16), .B(n38), .Z(\ab[34][3] ) );
  NR2 U602 ( .A(n15), .B(n38), .Z(\ab[34][2] ) );
  NR2 U603 ( .A(n5), .B(n38), .Z(\ab[34][21] ) );
  NR2 U604 ( .A(n6), .B(n38), .Z(\ab[34][20] ) );
  NR2 U605 ( .A(n14), .B(n38), .Z(\ab[34][1] ) );
  NR2 U606 ( .A(n7), .B(n38), .Z(\ab[34][19] ) );
  NR2 U607 ( .A(n8), .B(n38), .Z(\ab[34][18] ) );
  NR2 U608 ( .A(n9), .B(n38), .Z(\ab[34][17] ) );
  NR2 U609 ( .A(n10), .B(n38), .Z(\ab[34][16] ) );
  NR2 U610 ( .A(n11), .B(n38), .Z(\ab[34][15] ) );
  NR2 U611 ( .A(n4), .B(n38), .Z(\ab[34][14] ) );
  NR2 U612 ( .A(n12), .B(n38), .Z(\ab[34][13] ) );
  NR2 U613 ( .A(n25), .B(n38), .Z(\ab[34][12] ) );
  NR2 U614 ( .A(n24), .B(n38), .Z(\ab[34][11] ) );
  NR2 U615 ( .A(n23), .B(n38), .Z(\ab[34][10] ) );
  NR2 U616 ( .A(n13), .B(n38), .Z(\ab[34][0] ) );
  NR2 U617 ( .A(n22), .B(n39), .Z(\ab[33][9] ) );
  NR2 U618 ( .A(n21), .B(n39), .Z(\ab[33][8] ) );
  NR2 U619 ( .A(n20), .B(n39), .Z(\ab[33][7] ) );
  NR2 U620 ( .A(n19), .B(n39), .Z(\ab[33][6] ) );
  NR2 U621 ( .A(n18), .B(n39), .Z(\ab[33][5] ) );
  NR2 U622 ( .A(n17), .B(n39), .Z(\ab[33][4] ) );
  NR2 U623 ( .A(n16), .B(n39), .Z(\ab[33][3] ) );
  NR2 U624 ( .A(n15), .B(n39), .Z(\ab[33][2] ) );
  NR2 U625 ( .A(n5), .B(n39), .Z(\ab[33][21] ) );
  NR2 U626 ( .A(n6), .B(n39), .Z(\ab[33][20] ) );
  NR2 U627 ( .A(n14), .B(n39), .Z(\ab[33][1] ) );
  NR2 U628 ( .A(n7), .B(n39), .Z(\ab[33][19] ) );
  NR2 U629 ( .A(n8), .B(n39), .Z(\ab[33][18] ) );
  NR2 U630 ( .A(n9), .B(n39), .Z(\ab[33][17] ) );
  NR2 U631 ( .A(n10), .B(n39), .Z(\ab[33][16] ) );
  NR2 U632 ( .A(n11), .B(n39), .Z(\ab[33][15] ) );
  NR2 U633 ( .A(n4), .B(n39), .Z(\ab[33][14] ) );
  NR2 U634 ( .A(n12), .B(n39), .Z(\ab[33][13] ) );
  NR2 U635 ( .A(n25), .B(n39), .Z(\ab[33][12] ) );
  NR2 U636 ( .A(n24), .B(n39), .Z(\ab[33][11] ) );
  NR2 U637 ( .A(n23), .B(n39), .Z(\ab[33][10] ) );
  NR2 U638 ( .A(n13), .B(n39), .Z(\ab[33][0] ) );
  NR2 U639 ( .A(n22), .B(n40), .Z(\ab[32][9] ) );
  NR2 U640 ( .A(n21), .B(n40), .Z(\ab[32][8] ) );
  NR2 U641 ( .A(n20), .B(n40), .Z(\ab[32][7] ) );
  NR2 U642 ( .A(n19), .B(n40), .Z(\ab[32][6] ) );
  NR2 U643 ( .A(n18), .B(n40), .Z(\ab[32][5] ) );
  NR2 U644 ( .A(n17), .B(n40), .Z(\ab[32][4] ) );
  NR2 U645 ( .A(n16), .B(n40), .Z(\ab[32][3] ) );
  NR2 U646 ( .A(n15), .B(n40), .Z(\ab[32][2] ) );
  NR2 U647 ( .A(n5), .B(n40), .Z(\ab[32][21] ) );
  NR2 U648 ( .A(n6), .B(n40), .Z(\ab[32][20] ) );
  NR2 U649 ( .A(n14), .B(n40), .Z(\ab[32][1] ) );
  NR2 U650 ( .A(n7), .B(n40), .Z(\ab[32][19] ) );
  NR2 U651 ( .A(n8), .B(n40), .Z(\ab[32][18] ) );
  NR2 U652 ( .A(n9), .B(n40), .Z(\ab[32][17] ) );
  NR2 U653 ( .A(n10), .B(n40), .Z(\ab[32][16] ) );
  NR2 U654 ( .A(n11), .B(n40), .Z(\ab[32][15] ) );
  NR2 U655 ( .A(n4), .B(n40), .Z(\ab[32][14] ) );
  NR2 U656 ( .A(n12), .B(n40), .Z(\ab[32][13] ) );
  NR2 U657 ( .A(n25), .B(n40), .Z(\ab[32][12] ) );
  NR2 U658 ( .A(n24), .B(n40), .Z(\ab[32][11] ) );
  NR2 U659 ( .A(n23), .B(n40), .Z(\ab[32][10] ) );
  NR2 U660 ( .A(n13), .B(n40), .Z(\ab[32][0] ) );
  NR2 U661 ( .A(n22), .B(n41), .Z(\ab[31][9] ) );
  NR2 U662 ( .A(n21), .B(n41), .Z(\ab[31][8] ) );
  NR2 U663 ( .A(n20), .B(n41), .Z(\ab[31][7] ) );
  NR2 U664 ( .A(n19), .B(n41), .Z(\ab[31][6] ) );
  NR2 U665 ( .A(n18), .B(n41), .Z(\ab[31][5] ) );
  NR2 U666 ( .A(n17), .B(n41), .Z(\ab[31][4] ) );
  NR2 U667 ( .A(n16), .B(n41), .Z(\ab[31][3] ) );
  NR2 U668 ( .A(n15), .B(n41), .Z(\ab[31][2] ) );
  NR2 U669 ( .A(n5), .B(n41), .Z(\ab[31][21] ) );
  NR2 U670 ( .A(n6), .B(n41), .Z(\ab[31][20] ) );
  NR2 U671 ( .A(n14), .B(n41), .Z(\ab[31][1] ) );
  NR2 U672 ( .A(n7), .B(n41), .Z(\ab[31][19] ) );
  NR2 U673 ( .A(n8), .B(n41), .Z(\ab[31][18] ) );
  NR2 U674 ( .A(n9), .B(n41), .Z(\ab[31][17] ) );
  NR2 U675 ( .A(n10), .B(n41), .Z(\ab[31][16] ) );
  NR2 U676 ( .A(n11), .B(n41), .Z(\ab[31][15] ) );
  NR2 U677 ( .A(n4), .B(n41), .Z(\ab[31][14] ) );
  NR2 U678 ( .A(n12), .B(n41), .Z(\ab[31][13] ) );
  NR2 U679 ( .A(n25), .B(n41), .Z(\ab[31][12] ) );
  NR2 U680 ( .A(n24), .B(n41), .Z(\ab[31][11] ) );
  NR2 U681 ( .A(n23), .B(n41), .Z(\ab[31][10] ) );
  NR2 U682 ( .A(n13), .B(n41), .Z(\ab[31][0] ) );
  NR2 U683 ( .A(n22), .B(n42), .Z(\ab[30][9] ) );
  NR2 U684 ( .A(n21), .B(n42), .Z(\ab[30][8] ) );
  NR2 U685 ( .A(n20), .B(n42), .Z(\ab[30][7] ) );
  NR2 U686 ( .A(n19), .B(n42), .Z(\ab[30][6] ) );
  NR2 U687 ( .A(n18), .B(n42), .Z(\ab[30][5] ) );
  NR2 U688 ( .A(n17), .B(n42), .Z(\ab[30][4] ) );
  NR2 U689 ( .A(n16), .B(n42), .Z(\ab[30][3] ) );
  NR2 U690 ( .A(n15), .B(n42), .Z(\ab[30][2] ) );
  NR2 U691 ( .A(n5), .B(n42), .Z(\ab[30][21] ) );
  NR2 U692 ( .A(n6), .B(n42), .Z(\ab[30][20] ) );
  NR2 U693 ( .A(n14), .B(n42), .Z(\ab[30][1] ) );
  NR2 U694 ( .A(n7), .B(n42), .Z(\ab[30][19] ) );
  NR2 U695 ( .A(n8), .B(n42), .Z(\ab[30][18] ) );
  NR2 U696 ( .A(n9), .B(n42), .Z(\ab[30][17] ) );
  NR2 U697 ( .A(n10), .B(n42), .Z(\ab[30][16] ) );
  NR2 U698 ( .A(n11), .B(n42), .Z(\ab[30][15] ) );
  NR2 U699 ( .A(n4), .B(n42), .Z(\ab[30][14] ) );
  NR2 U700 ( .A(n12), .B(n42), .Z(\ab[30][13] ) );
  NR2 U701 ( .A(n25), .B(n42), .Z(\ab[30][12] ) );
  NR2 U702 ( .A(n24), .B(n42), .Z(\ab[30][11] ) );
  NR2 U703 ( .A(n23), .B(n42), .Z(\ab[30][10] ) );
  NR2 U704 ( .A(n13), .B(n42), .Z(\ab[30][0] ) );
  NR2 U705 ( .A(n22), .B(n70), .Z(\ab[2][9] ) );
  NR2 U706 ( .A(n21), .B(n70), .Z(\ab[2][8] ) );
  NR2 U707 ( .A(n20), .B(n70), .Z(\ab[2][7] ) );
  NR2 U708 ( .A(n19), .B(n70), .Z(\ab[2][6] ) );
  NR2 U709 ( .A(n18), .B(n70), .Z(\ab[2][5] ) );
  NR2 U710 ( .A(n17), .B(n70), .Z(\ab[2][4] ) );
  NR2 U711 ( .A(n16), .B(n70), .Z(\ab[2][3] ) );
  NR2 U712 ( .A(n15), .B(n70), .Z(\ab[2][2] ) );
  NR2 U713 ( .A(n5), .B(n70), .Z(\ab[2][21] ) );
  NR2 U714 ( .A(n6), .B(n70), .Z(\ab[2][20] ) );
  NR2 U715 ( .A(n14), .B(n70), .Z(\ab[2][1] ) );
  NR2 U716 ( .A(n7), .B(n70), .Z(\ab[2][19] ) );
  NR2 U717 ( .A(n8), .B(n70), .Z(\ab[2][18] ) );
  NR2 U718 ( .A(n9), .B(n70), .Z(\ab[2][17] ) );
  NR2 U719 ( .A(n10), .B(n70), .Z(\ab[2][16] ) );
  NR2 U720 ( .A(n11), .B(n70), .Z(\ab[2][15] ) );
  NR2 U721 ( .A(n4), .B(n70), .Z(\ab[2][14] ) );
  NR2 U722 ( .A(n12), .B(n70), .Z(\ab[2][13] ) );
  NR2 U723 ( .A(n25), .B(n70), .Z(\ab[2][12] ) );
  NR2 U724 ( .A(n24), .B(n70), .Z(\ab[2][11] ) );
  NR2 U725 ( .A(n23), .B(n70), .Z(\ab[2][10] ) );
  NR2 U726 ( .A(n13), .B(n70), .Z(\ab[2][0] ) );
  NR2 U727 ( .A(n22), .B(n43), .Z(\ab[29][9] ) );
  NR2 U728 ( .A(n21), .B(n43), .Z(\ab[29][8] ) );
  NR2 U729 ( .A(n20), .B(n43), .Z(\ab[29][7] ) );
  NR2 U730 ( .A(n19), .B(n43), .Z(\ab[29][6] ) );
  NR2 U731 ( .A(n18), .B(n43), .Z(\ab[29][5] ) );
  NR2 U732 ( .A(n17), .B(n43), .Z(\ab[29][4] ) );
  NR2 U733 ( .A(n16), .B(n43), .Z(\ab[29][3] ) );
  NR2 U734 ( .A(n15), .B(n43), .Z(\ab[29][2] ) );
  NR2 U735 ( .A(n5), .B(n43), .Z(\ab[29][21] ) );
  NR2 U736 ( .A(n6), .B(n43), .Z(\ab[29][20] ) );
  NR2 U737 ( .A(n14), .B(n43), .Z(\ab[29][1] ) );
  NR2 U738 ( .A(n7), .B(n43), .Z(\ab[29][19] ) );
  NR2 U739 ( .A(n8), .B(n43), .Z(\ab[29][18] ) );
  NR2 U740 ( .A(n9), .B(n43), .Z(\ab[29][17] ) );
  NR2 U741 ( .A(n10), .B(n43), .Z(\ab[29][16] ) );
  NR2 U742 ( .A(n11), .B(n43), .Z(\ab[29][15] ) );
  NR2 U743 ( .A(n4), .B(n43), .Z(\ab[29][14] ) );
  NR2 U744 ( .A(n12), .B(n43), .Z(\ab[29][13] ) );
  NR2 U745 ( .A(n25), .B(n43), .Z(\ab[29][12] ) );
  NR2 U746 ( .A(n24), .B(n43), .Z(\ab[29][11] ) );
  NR2 U747 ( .A(n23), .B(n43), .Z(\ab[29][10] ) );
  NR2 U748 ( .A(n13), .B(n43), .Z(\ab[29][0] ) );
  NR2 U749 ( .A(n22), .B(n44), .Z(\ab[28][9] ) );
  NR2 U750 ( .A(n21), .B(n44), .Z(\ab[28][8] ) );
  NR2 U751 ( .A(n20), .B(n44), .Z(\ab[28][7] ) );
  NR2 U752 ( .A(n19), .B(n44), .Z(\ab[28][6] ) );
  NR2 U753 ( .A(n18), .B(n44), .Z(\ab[28][5] ) );
  NR2 U754 ( .A(n17), .B(n44), .Z(\ab[28][4] ) );
  NR2 U755 ( .A(n16), .B(n44), .Z(\ab[28][3] ) );
  NR2 U756 ( .A(n15), .B(n44), .Z(\ab[28][2] ) );
  NR2 U757 ( .A(n5), .B(n44), .Z(\ab[28][21] ) );
  NR2 U758 ( .A(n6), .B(n44), .Z(\ab[28][20] ) );
  NR2 U759 ( .A(n14), .B(n44), .Z(\ab[28][1] ) );
  NR2 U760 ( .A(n7), .B(n44), .Z(\ab[28][19] ) );
  NR2 U761 ( .A(n8), .B(n44), .Z(\ab[28][18] ) );
  NR2 U762 ( .A(n9), .B(n44), .Z(\ab[28][17] ) );
  NR2 U763 ( .A(n10), .B(n44), .Z(\ab[28][16] ) );
  NR2 U764 ( .A(n11), .B(n44), .Z(\ab[28][15] ) );
  NR2 U765 ( .A(n4), .B(n44), .Z(\ab[28][14] ) );
  NR2 U766 ( .A(n12), .B(n44), .Z(\ab[28][13] ) );
  NR2 U767 ( .A(n25), .B(n44), .Z(\ab[28][12] ) );
  NR2 U768 ( .A(n24), .B(n44), .Z(\ab[28][11] ) );
  NR2 U769 ( .A(n23), .B(n44), .Z(\ab[28][10] ) );
  NR2 U770 ( .A(n13), .B(n44), .Z(\ab[28][0] ) );
  NR2 U771 ( .A(n22), .B(n45), .Z(\ab[27][9] ) );
  NR2 U772 ( .A(n21), .B(n45), .Z(\ab[27][8] ) );
  NR2 U773 ( .A(n20), .B(n45), .Z(\ab[27][7] ) );
  NR2 U774 ( .A(n19), .B(n45), .Z(\ab[27][6] ) );
  NR2 U775 ( .A(n18), .B(n45), .Z(\ab[27][5] ) );
  NR2 U776 ( .A(n17), .B(n45), .Z(\ab[27][4] ) );
  NR2 U777 ( .A(n16), .B(n45), .Z(\ab[27][3] ) );
  NR2 U778 ( .A(n15), .B(n45), .Z(\ab[27][2] ) );
  NR2 U779 ( .A(n5), .B(n45), .Z(\ab[27][21] ) );
  NR2 U780 ( .A(n6), .B(n45), .Z(\ab[27][20] ) );
  NR2 U781 ( .A(n14), .B(n45), .Z(\ab[27][1] ) );
  NR2 U782 ( .A(n7), .B(n45), .Z(\ab[27][19] ) );
  NR2 U783 ( .A(n8), .B(n45), .Z(\ab[27][18] ) );
  NR2 U784 ( .A(n9), .B(n45), .Z(\ab[27][17] ) );
  NR2 U785 ( .A(n10), .B(n45), .Z(\ab[27][16] ) );
  NR2 U786 ( .A(n11), .B(n45), .Z(\ab[27][15] ) );
  NR2 U787 ( .A(n4), .B(n45), .Z(\ab[27][14] ) );
  NR2 U788 ( .A(n12), .B(n45), .Z(\ab[27][13] ) );
  NR2 U789 ( .A(n25), .B(n45), .Z(\ab[27][12] ) );
  NR2 U790 ( .A(n24), .B(n45), .Z(\ab[27][11] ) );
  NR2 U791 ( .A(n23), .B(n45), .Z(\ab[27][10] ) );
  NR2 U792 ( .A(n13), .B(n45), .Z(\ab[27][0] ) );
  NR2 U793 ( .A(n22), .B(n46), .Z(\ab[26][9] ) );
  NR2 U794 ( .A(n21), .B(n46), .Z(\ab[26][8] ) );
  NR2 U795 ( .A(n20), .B(n46), .Z(\ab[26][7] ) );
  NR2 U796 ( .A(n19), .B(n46), .Z(\ab[26][6] ) );
  NR2 U797 ( .A(n18), .B(n46), .Z(\ab[26][5] ) );
  NR2 U798 ( .A(n17), .B(n46), .Z(\ab[26][4] ) );
  NR2 U799 ( .A(n16), .B(n46), .Z(\ab[26][3] ) );
  NR2 U800 ( .A(n15), .B(n46), .Z(\ab[26][2] ) );
  NR2 U801 ( .A(n5), .B(n46), .Z(\ab[26][21] ) );
  NR2 U802 ( .A(n6), .B(n46), .Z(\ab[26][20] ) );
  NR2 U803 ( .A(n14), .B(n46), .Z(\ab[26][1] ) );
  NR2 U804 ( .A(n7), .B(n46), .Z(\ab[26][19] ) );
  NR2 U805 ( .A(n8), .B(n46), .Z(\ab[26][18] ) );
  NR2 U806 ( .A(n9), .B(n46), .Z(\ab[26][17] ) );
  NR2 U807 ( .A(n10), .B(n46), .Z(\ab[26][16] ) );
  NR2 U808 ( .A(n11), .B(n46), .Z(\ab[26][15] ) );
  NR2 U809 ( .A(n4), .B(n46), .Z(\ab[26][14] ) );
  NR2 U810 ( .A(n12), .B(n46), .Z(\ab[26][13] ) );
  NR2 U811 ( .A(n25), .B(n46), .Z(\ab[26][12] ) );
  NR2 U812 ( .A(n24), .B(n46), .Z(\ab[26][11] ) );
  NR2 U813 ( .A(n23), .B(n46), .Z(\ab[26][10] ) );
  NR2 U814 ( .A(n13), .B(n46), .Z(\ab[26][0] ) );
  NR2 U815 ( .A(n22), .B(n47), .Z(\ab[25][9] ) );
  NR2 U816 ( .A(n21), .B(n47), .Z(\ab[25][8] ) );
  NR2 U817 ( .A(n20), .B(n47), .Z(\ab[25][7] ) );
  NR2 U818 ( .A(n19), .B(n47), .Z(\ab[25][6] ) );
  NR2 U819 ( .A(n18), .B(n47), .Z(\ab[25][5] ) );
  NR2 U820 ( .A(n17), .B(n47), .Z(\ab[25][4] ) );
  NR2 U821 ( .A(n16), .B(n47), .Z(\ab[25][3] ) );
  NR2 U822 ( .A(n15), .B(n47), .Z(\ab[25][2] ) );
  NR2 U823 ( .A(n5), .B(n47), .Z(\ab[25][21] ) );
  NR2 U824 ( .A(n6), .B(n47), .Z(\ab[25][20] ) );
  NR2 U825 ( .A(n14), .B(n47), .Z(\ab[25][1] ) );
  NR2 U826 ( .A(n7), .B(n47), .Z(\ab[25][19] ) );
  NR2 U827 ( .A(n8), .B(n47), .Z(\ab[25][18] ) );
  NR2 U828 ( .A(n9), .B(n47), .Z(\ab[25][17] ) );
  NR2 U829 ( .A(n10), .B(n47), .Z(\ab[25][16] ) );
  NR2 U830 ( .A(n11), .B(n47), .Z(\ab[25][15] ) );
  NR2 U831 ( .A(n4), .B(n47), .Z(\ab[25][14] ) );
  NR2 U832 ( .A(n12), .B(n47), .Z(\ab[25][13] ) );
  NR2 U833 ( .A(n25), .B(n47), .Z(\ab[25][12] ) );
  NR2 U834 ( .A(n24), .B(n47), .Z(\ab[25][11] ) );
  NR2 U835 ( .A(n23), .B(n47), .Z(\ab[25][10] ) );
  NR2 U836 ( .A(n13), .B(n47), .Z(\ab[25][0] ) );
  NR2 U837 ( .A(n22), .B(n48), .Z(\ab[24][9] ) );
  NR2 U838 ( .A(n21), .B(n48), .Z(\ab[24][8] ) );
  NR2 U839 ( .A(n20), .B(n48), .Z(\ab[24][7] ) );
  NR2 U840 ( .A(n19), .B(n48), .Z(\ab[24][6] ) );
  NR2 U841 ( .A(n18), .B(n48), .Z(\ab[24][5] ) );
  NR2 U842 ( .A(n17), .B(n48), .Z(\ab[24][4] ) );
  NR2 U843 ( .A(n16), .B(n48), .Z(\ab[24][3] ) );
  NR2 U844 ( .A(n15), .B(n48), .Z(\ab[24][2] ) );
  NR2 U845 ( .A(n5), .B(n48), .Z(\ab[24][21] ) );
  NR2 U846 ( .A(n6), .B(n48), .Z(\ab[24][20] ) );
  NR2 U847 ( .A(n14), .B(n48), .Z(\ab[24][1] ) );
  NR2 U848 ( .A(n7), .B(n48), .Z(\ab[24][19] ) );
  NR2 U849 ( .A(n8), .B(n48), .Z(\ab[24][18] ) );
  NR2 U850 ( .A(n9), .B(n48), .Z(\ab[24][17] ) );
  NR2 U851 ( .A(n10), .B(n48), .Z(\ab[24][16] ) );
  NR2 U852 ( .A(n11), .B(n48), .Z(\ab[24][15] ) );
  NR2 U853 ( .A(n4), .B(n48), .Z(\ab[24][14] ) );
  NR2 U854 ( .A(n12), .B(n48), .Z(\ab[24][13] ) );
  NR2 U855 ( .A(n25), .B(n48), .Z(\ab[24][12] ) );
  NR2 U856 ( .A(n24), .B(n48), .Z(\ab[24][11] ) );
  NR2 U857 ( .A(n23), .B(n48), .Z(\ab[24][10] ) );
  NR2 U858 ( .A(n13), .B(n48), .Z(\ab[24][0] ) );
  NR2 U859 ( .A(n22), .B(n49), .Z(\ab[23][9] ) );
  NR2 U860 ( .A(n21), .B(n49), .Z(\ab[23][8] ) );
  NR2 U861 ( .A(n20), .B(n49), .Z(\ab[23][7] ) );
  NR2 U862 ( .A(n19), .B(n49), .Z(\ab[23][6] ) );
  NR2 U863 ( .A(n18), .B(n49), .Z(\ab[23][5] ) );
  NR2 U864 ( .A(n17), .B(n49), .Z(\ab[23][4] ) );
  NR2 U865 ( .A(n16), .B(n49), .Z(\ab[23][3] ) );
  NR2 U866 ( .A(n15), .B(n49), .Z(\ab[23][2] ) );
  NR2 U867 ( .A(n5), .B(n49), .Z(\ab[23][21] ) );
  NR2 U868 ( .A(n6), .B(n49), .Z(\ab[23][20] ) );
  NR2 U869 ( .A(n14), .B(n49), .Z(\ab[23][1] ) );
  NR2 U870 ( .A(n7), .B(n49), .Z(\ab[23][19] ) );
  NR2 U871 ( .A(n8), .B(n49), .Z(\ab[23][18] ) );
  NR2 U872 ( .A(n9), .B(n49), .Z(\ab[23][17] ) );
  NR2 U873 ( .A(n10), .B(n49), .Z(\ab[23][16] ) );
  NR2 U874 ( .A(n11), .B(n49), .Z(\ab[23][15] ) );
  NR2 U875 ( .A(n4), .B(n49), .Z(\ab[23][14] ) );
  NR2 U876 ( .A(n12), .B(n49), .Z(\ab[23][13] ) );
  NR2 U877 ( .A(n25), .B(n49), .Z(\ab[23][12] ) );
  NR2 U878 ( .A(n24), .B(n49), .Z(\ab[23][11] ) );
  NR2 U879 ( .A(n23), .B(n49), .Z(\ab[23][10] ) );
  NR2 U880 ( .A(n13), .B(n49), .Z(\ab[23][0] ) );
  NR2 U881 ( .A(n22), .B(n50), .Z(\ab[22][9] ) );
  NR2 U882 ( .A(n21), .B(n50), .Z(\ab[22][8] ) );
  NR2 U883 ( .A(n20), .B(n50), .Z(\ab[22][7] ) );
  NR2 U884 ( .A(n19), .B(n50), .Z(\ab[22][6] ) );
  NR2 U885 ( .A(n18), .B(n50), .Z(\ab[22][5] ) );
  NR2 U886 ( .A(n17), .B(n50), .Z(\ab[22][4] ) );
  NR2 U887 ( .A(n16), .B(n50), .Z(\ab[22][3] ) );
  NR2 U888 ( .A(n15), .B(n50), .Z(\ab[22][2] ) );
  NR2 U889 ( .A(n5), .B(n50), .Z(\ab[22][21] ) );
  NR2 U890 ( .A(n6), .B(n50), .Z(\ab[22][20] ) );
  NR2 U891 ( .A(n14), .B(n50), .Z(\ab[22][1] ) );
  NR2 U892 ( .A(n7), .B(n50), .Z(\ab[22][19] ) );
  NR2 U893 ( .A(n8), .B(n50), .Z(\ab[22][18] ) );
  NR2 U894 ( .A(n9), .B(n50), .Z(\ab[22][17] ) );
  NR2 U895 ( .A(n10), .B(n50), .Z(\ab[22][16] ) );
  NR2 U896 ( .A(n11), .B(n50), .Z(\ab[22][15] ) );
  NR2 U897 ( .A(n4), .B(n50), .Z(\ab[22][14] ) );
  NR2 U898 ( .A(n12), .B(n50), .Z(\ab[22][13] ) );
  NR2 U899 ( .A(n25), .B(n50), .Z(\ab[22][12] ) );
  NR2 U900 ( .A(n24), .B(n50), .Z(\ab[22][11] ) );
  NR2 U901 ( .A(n23), .B(n50), .Z(\ab[22][10] ) );
  NR2 U902 ( .A(n13), .B(n50), .Z(\ab[22][0] ) );
  NR2 U903 ( .A(n22), .B(n51), .Z(\ab[21][9] ) );
  NR2 U904 ( .A(n21), .B(n51), .Z(\ab[21][8] ) );
  NR2 U905 ( .A(n20), .B(n51), .Z(\ab[21][7] ) );
  NR2 U906 ( .A(n19), .B(n51), .Z(\ab[21][6] ) );
  NR2 U907 ( .A(n18), .B(n51), .Z(\ab[21][5] ) );
  NR2 U908 ( .A(n17), .B(n51), .Z(\ab[21][4] ) );
  NR2 U909 ( .A(n16), .B(n51), .Z(\ab[21][3] ) );
  NR2 U910 ( .A(n15), .B(n51), .Z(\ab[21][2] ) );
  NR2 U911 ( .A(n5), .B(n51), .Z(\ab[21][21] ) );
  NR2 U912 ( .A(n6), .B(n51), .Z(\ab[21][20] ) );
  NR2 U913 ( .A(n14), .B(n51), .Z(\ab[21][1] ) );
  NR2 U914 ( .A(n7), .B(n51), .Z(\ab[21][19] ) );
  NR2 U915 ( .A(n8), .B(n51), .Z(\ab[21][18] ) );
  NR2 U916 ( .A(n9), .B(n51), .Z(\ab[21][17] ) );
  NR2 U917 ( .A(n10), .B(n51), .Z(\ab[21][16] ) );
  NR2 U918 ( .A(n11), .B(n51), .Z(\ab[21][15] ) );
  NR2 U919 ( .A(n4), .B(n51), .Z(\ab[21][14] ) );
  NR2 U920 ( .A(n12), .B(n51), .Z(\ab[21][13] ) );
  NR2 U921 ( .A(n25), .B(n51), .Z(\ab[21][12] ) );
  NR2 U922 ( .A(n24), .B(n51), .Z(\ab[21][11] ) );
  NR2 U923 ( .A(n23), .B(n51), .Z(\ab[21][10] ) );
  NR2 U924 ( .A(n13), .B(n51), .Z(\ab[21][0] ) );
  NR2 U925 ( .A(n22), .B(n52), .Z(\ab[20][9] ) );
  NR2 U926 ( .A(n21), .B(n52), .Z(\ab[20][8] ) );
  NR2 U927 ( .A(n20), .B(n52), .Z(\ab[20][7] ) );
  NR2 U928 ( .A(n19), .B(n52), .Z(\ab[20][6] ) );
  NR2 U929 ( .A(n18), .B(n52), .Z(\ab[20][5] ) );
  NR2 U930 ( .A(n17), .B(n52), .Z(\ab[20][4] ) );
  NR2 U931 ( .A(n16), .B(n52), .Z(\ab[20][3] ) );
  NR2 U932 ( .A(n15), .B(n52), .Z(\ab[20][2] ) );
  NR2 U933 ( .A(n5), .B(n52), .Z(\ab[20][21] ) );
  NR2 U934 ( .A(n6), .B(n52), .Z(\ab[20][20] ) );
  NR2 U935 ( .A(n14), .B(n52), .Z(\ab[20][1] ) );
  NR2 U936 ( .A(n7), .B(n52), .Z(\ab[20][19] ) );
  NR2 U937 ( .A(n8), .B(n52), .Z(\ab[20][18] ) );
  NR2 U938 ( .A(n9), .B(n52), .Z(\ab[20][17] ) );
  NR2 U939 ( .A(n10), .B(n52), .Z(\ab[20][16] ) );
  NR2 U940 ( .A(n11), .B(n52), .Z(\ab[20][15] ) );
  NR2 U941 ( .A(n4), .B(n52), .Z(\ab[20][14] ) );
  NR2 U942 ( .A(n12), .B(n52), .Z(\ab[20][13] ) );
  NR2 U943 ( .A(n25), .B(n52), .Z(\ab[20][12] ) );
  NR2 U944 ( .A(n24), .B(n52), .Z(\ab[20][11] ) );
  NR2 U945 ( .A(n23), .B(n52), .Z(\ab[20][10] ) );
  NR2 U946 ( .A(n13), .B(n52), .Z(\ab[20][0] ) );
  NR2 U947 ( .A(n22), .B(n71), .Z(\ab[1][9] ) );
  NR2 U948 ( .A(n21), .B(n71), .Z(\ab[1][8] ) );
  NR2 U949 ( .A(n20), .B(n71), .Z(\ab[1][7] ) );
  NR2 U950 ( .A(n19), .B(n71), .Z(\ab[1][6] ) );
  NR2 U951 ( .A(n18), .B(n71), .Z(\ab[1][5] ) );
  NR2 U952 ( .A(n17), .B(n71), .Z(\ab[1][4] ) );
  NR2 U953 ( .A(n16), .B(n71), .Z(\ab[1][3] ) );
  NR2 U954 ( .A(n15), .B(n71), .Z(\ab[1][2] ) );
  NR2 U955 ( .A(n5), .B(n71), .Z(\ab[1][21] ) );
  NR2 U956 ( .A(n6), .B(n71), .Z(\ab[1][20] ) );
  NR2 U957 ( .A(n7), .B(n71), .Z(\ab[1][19] ) );
  NR2 U958 ( .A(n8), .B(n71), .Z(\ab[1][18] ) );
  NR2 U959 ( .A(n9), .B(n71), .Z(\ab[1][17] ) );
  NR2 U960 ( .A(n10), .B(n71), .Z(\ab[1][16] ) );
  NR2 U961 ( .A(n11), .B(n71), .Z(\ab[1][15] ) );
  NR2 U962 ( .A(n4), .B(n71), .Z(\ab[1][14] ) );
  NR2 U963 ( .A(n12), .B(n71), .Z(\ab[1][13] ) );
  NR2 U964 ( .A(n25), .B(n71), .Z(\ab[1][12] ) );
  NR2 U965 ( .A(n24), .B(n71), .Z(\ab[1][11] ) );
  NR2 U966 ( .A(n23), .B(n71), .Z(\ab[1][10] ) );
  NR2 U967 ( .A(n22), .B(n53), .Z(\ab[19][9] ) );
  NR2 U968 ( .A(n21), .B(n53), .Z(\ab[19][8] ) );
  NR2 U969 ( .A(n20), .B(n53), .Z(\ab[19][7] ) );
  NR2 U970 ( .A(n19), .B(n53), .Z(\ab[19][6] ) );
  NR2 U971 ( .A(n18), .B(n53), .Z(\ab[19][5] ) );
  NR2 U972 ( .A(n17), .B(n53), .Z(\ab[19][4] ) );
  NR2 U973 ( .A(n16), .B(n53), .Z(\ab[19][3] ) );
  NR2 U974 ( .A(n15), .B(n53), .Z(\ab[19][2] ) );
  NR2 U975 ( .A(n5), .B(n53), .Z(\ab[19][21] ) );
  NR2 U976 ( .A(n6), .B(n53), .Z(\ab[19][20] ) );
  NR2 U977 ( .A(n14), .B(n53), .Z(\ab[19][1] ) );
  NR2 U978 ( .A(n7), .B(n53), .Z(\ab[19][19] ) );
  NR2 U979 ( .A(n8), .B(n53), .Z(\ab[19][18] ) );
  NR2 U980 ( .A(n9), .B(n53), .Z(\ab[19][17] ) );
  NR2 U981 ( .A(n10), .B(n53), .Z(\ab[19][16] ) );
  NR2 U982 ( .A(n11), .B(n53), .Z(\ab[19][15] ) );
  NR2 U983 ( .A(n4), .B(n53), .Z(\ab[19][14] ) );
  NR2 U984 ( .A(n12), .B(n53), .Z(\ab[19][13] ) );
  NR2 U985 ( .A(n25), .B(n53), .Z(\ab[19][12] ) );
  NR2 U986 ( .A(n24), .B(n53), .Z(\ab[19][11] ) );
  NR2 U987 ( .A(n23), .B(n53), .Z(\ab[19][10] ) );
  NR2 U988 ( .A(n13), .B(n53), .Z(\ab[19][0] ) );
  NR2 U989 ( .A(n22), .B(n54), .Z(\ab[18][9] ) );
  NR2 U990 ( .A(n21), .B(n54), .Z(\ab[18][8] ) );
  NR2 U991 ( .A(n20), .B(n54), .Z(\ab[18][7] ) );
  NR2 U992 ( .A(n19), .B(n54), .Z(\ab[18][6] ) );
  NR2 U993 ( .A(n18), .B(n54), .Z(\ab[18][5] ) );
  NR2 U994 ( .A(n17), .B(n54), .Z(\ab[18][4] ) );
  NR2 U995 ( .A(n16), .B(n54), .Z(\ab[18][3] ) );
  NR2 U996 ( .A(n15), .B(n54), .Z(\ab[18][2] ) );
  NR2 U997 ( .A(n5), .B(n54), .Z(\ab[18][21] ) );
  NR2 U998 ( .A(n6), .B(n54), .Z(\ab[18][20] ) );
  NR2 U999 ( .A(n14), .B(n54), .Z(\ab[18][1] ) );
  NR2 U1000 ( .A(n7), .B(n54), .Z(\ab[18][19] ) );
  NR2 U1001 ( .A(n8), .B(n54), .Z(\ab[18][18] ) );
  NR2 U1002 ( .A(n9), .B(n54), .Z(\ab[18][17] ) );
  NR2 U1003 ( .A(n10), .B(n54), .Z(\ab[18][16] ) );
  NR2 U1004 ( .A(n11), .B(n54), .Z(\ab[18][15] ) );
  NR2 U1005 ( .A(n4), .B(n54), .Z(\ab[18][14] ) );
  NR2 U1006 ( .A(n12), .B(n54), .Z(\ab[18][13] ) );
  NR2 U1007 ( .A(n25), .B(n54), .Z(\ab[18][12] ) );
  NR2 U1008 ( .A(n24), .B(n54), .Z(\ab[18][11] ) );
  NR2 U1009 ( .A(n23), .B(n54), .Z(\ab[18][10] ) );
  NR2 U1010 ( .A(n13), .B(n54), .Z(\ab[18][0] ) );
  NR2 U1011 ( .A(n22), .B(n55), .Z(\ab[17][9] ) );
  NR2 U1012 ( .A(n21), .B(n55), .Z(\ab[17][8] ) );
  NR2 U1013 ( .A(n20), .B(n55), .Z(\ab[17][7] ) );
  NR2 U1014 ( .A(n19), .B(n55), .Z(\ab[17][6] ) );
  NR2 U1015 ( .A(n18), .B(n55), .Z(\ab[17][5] ) );
  NR2 U1016 ( .A(n17), .B(n55), .Z(\ab[17][4] ) );
  NR2 U1017 ( .A(n16), .B(n55), .Z(\ab[17][3] ) );
  NR2 U1018 ( .A(n15), .B(n55), .Z(\ab[17][2] ) );
  NR2 U1019 ( .A(n5), .B(n55), .Z(\ab[17][21] ) );
  NR2 U1020 ( .A(n6), .B(n55), .Z(\ab[17][20] ) );
  NR2 U1021 ( .A(n14), .B(n55), .Z(\ab[17][1] ) );
  NR2 U1022 ( .A(n7), .B(n55), .Z(\ab[17][19] ) );
  NR2 U1023 ( .A(n8), .B(n55), .Z(\ab[17][18] ) );
  NR2 U1024 ( .A(n9), .B(n55), .Z(\ab[17][17] ) );
  NR2 U1025 ( .A(n10), .B(n55), .Z(\ab[17][16] ) );
  NR2 U1026 ( .A(n11), .B(n55), .Z(\ab[17][15] ) );
  NR2 U1027 ( .A(n4), .B(n55), .Z(\ab[17][14] ) );
  NR2 U1028 ( .A(n12), .B(n55), .Z(\ab[17][13] ) );
  NR2 U1029 ( .A(n25), .B(n55), .Z(\ab[17][12] ) );
  NR2 U1030 ( .A(n24), .B(n55), .Z(\ab[17][11] ) );
  NR2 U1031 ( .A(n23), .B(n55), .Z(\ab[17][10] ) );
  NR2 U1032 ( .A(n13), .B(n55), .Z(\ab[17][0] ) );
  NR2 U1033 ( .A(n22), .B(n56), .Z(\ab[16][9] ) );
  NR2 U1034 ( .A(n21), .B(n56), .Z(\ab[16][8] ) );
  NR2 U1035 ( .A(n20), .B(n56), .Z(\ab[16][7] ) );
  NR2 U1036 ( .A(n19), .B(n56), .Z(\ab[16][6] ) );
  NR2 U1037 ( .A(n18), .B(n56), .Z(\ab[16][5] ) );
  NR2 U1038 ( .A(n17), .B(n56), .Z(\ab[16][4] ) );
  NR2 U1039 ( .A(n16), .B(n56), .Z(\ab[16][3] ) );
  NR2 U1040 ( .A(n15), .B(n56), .Z(\ab[16][2] ) );
  NR2 U1041 ( .A(n5), .B(n56), .Z(\ab[16][21] ) );
  NR2 U1042 ( .A(n6), .B(n56), .Z(\ab[16][20] ) );
  NR2 U1043 ( .A(n14), .B(n56), .Z(\ab[16][1] ) );
  NR2 U1044 ( .A(n7), .B(n56), .Z(\ab[16][19] ) );
  NR2 U1045 ( .A(n8), .B(n56), .Z(\ab[16][18] ) );
  NR2 U1046 ( .A(n9), .B(n56), .Z(\ab[16][17] ) );
  NR2 U1047 ( .A(n10), .B(n56), .Z(\ab[16][16] ) );
  NR2 U1048 ( .A(n11), .B(n56), .Z(\ab[16][15] ) );
  NR2 U1049 ( .A(n4), .B(n56), .Z(\ab[16][14] ) );
  NR2 U1050 ( .A(n12), .B(n56), .Z(\ab[16][13] ) );
  NR2 U1051 ( .A(n25), .B(n56), .Z(\ab[16][12] ) );
  NR2 U1052 ( .A(n24), .B(n56), .Z(\ab[16][11] ) );
  NR2 U1053 ( .A(n23), .B(n56), .Z(\ab[16][10] ) );
  NR2 U1054 ( .A(n13), .B(n56), .Z(\ab[16][0] ) );
  NR2 U1055 ( .A(n22), .B(n57), .Z(\ab[15][9] ) );
  NR2 U1056 ( .A(n21), .B(n57), .Z(\ab[15][8] ) );
  NR2 U1057 ( .A(n20), .B(n57), .Z(\ab[15][7] ) );
  NR2 U1058 ( .A(n19), .B(n57), .Z(\ab[15][6] ) );
  NR2 U1059 ( .A(n18), .B(n57), .Z(\ab[15][5] ) );
  NR2 U1060 ( .A(n17), .B(n57), .Z(\ab[15][4] ) );
  NR2 U1061 ( .A(n16), .B(n57), .Z(\ab[15][3] ) );
  NR2 U1062 ( .A(n15), .B(n57), .Z(\ab[15][2] ) );
  NR2 U1063 ( .A(n5), .B(n57), .Z(\ab[15][21] ) );
  NR2 U1064 ( .A(n6), .B(n57), .Z(\ab[15][20] ) );
  NR2 U1065 ( .A(n14), .B(n57), .Z(\ab[15][1] ) );
  NR2 U1066 ( .A(n7), .B(n57), .Z(\ab[15][19] ) );
  NR2 U1067 ( .A(n8), .B(n57), .Z(\ab[15][18] ) );
  NR2 U1068 ( .A(n9), .B(n57), .Z(\ab[15][17] ) );
  NR2 U1069 ( .A(n10), .B(n57), .Z(\ab[15][16] ) );
  NR2 U1070 ( .A(n11), .B(n57), .Z(\ab[15][15] ) );
  NR2 U1071 ( .A(n4), .B(n57), .Z(\ab[15][14] ) );
  NR2 U1072 ( .A(n12), .B(n57), .Z(\ab[15][13] ) );
  NR2 U1073 ( .A(n25), .B(n57), .Z(\ab[15][12] ) );
  NR2 U1074 ( .A(n24), .B(n57), .Z(\ab[15][11] ) );
  NR2 U1075 ( .A(n23), .B(n57), .Z(\ab[15][10] ) );
  NR2 U1076 ( .A(n13), .B(n57), .Z(\ab[15][0] ) );
  NR2 U1077 ( .A(n22), .B(n58), .Z(\ab[14][9] ) );
  NR2 U1078 ( .A(n21), .B(n58), .Z(\ab[14][8] ) );
  NR2 U1079 ( .A(n20), .B(n58), .Z(\ab[14][7] ) );
  NR2 U1080 ( .A(n19), .B(n58), .Z(\ab[14][6] ) );
  NR2 U1081 ( .A(n18), .B(n58), .Z(\ab[14][5] ) );
  NR2 U1082 ( .A(n17), .B(n58), .Z(\ab[14][4] ) );
  NR2 U1083 ( .A(n16), .B(n58), .Z(\ab[14][3] ) );
  NR2 U1084 ( .A(n15), .B(n58), .Z(\ab[14][2] ) );
  NR2 U1085 ( .A(n5), .B(n58), .Z(\ab[14][21] ) );
  NR2 U1086 ( .A(n6), .B(n58), .Z(\ab[14][20] ) );
  NR2 U1087 ( .A(n14), .B(n58), .Z(\ab[14][1] ) );
  NR2 U1088 ( .A(n7), .B(n58), .Z(\ab[14][19] ) );
  NR2 U1089 ( .A(n8), .B(n58), .Z(\ab[14][18] ) );
  NR2 U1090 ( .A(n9), .B(n58), .Z(\ab[14][17] ) );
  NR2 U1091 ( .A(n10), .B(n58), .Z(\ab[14][16] ) );
  NR2 U1092 ( .A(n11), .B(n58), .Z(\ab[14][15] ) );
  NR2 U1093 ( .A(n4), .B(n58), .Z(\ab[14][14] ) );
  NR2 U1094 ( .A(n12), .B(n58), .Z(\ab[14][13] ) );
  NR2 U1095 ( .A(n25), .B(n58), .Z(\ab[14][12] ) );
  NR2 U1096 ( .A(n24), .B(n58), .Z(\ab[14][11] ) );
  NR2 U1097 ( .A(n23), .B(n58), .Z(\ab[14][10] ) );
  NR2 U1098 ( .A(n13), .B(n58), .Z(\ab[14][0] ) );
  NR2 U1099 ( .A(n22), .B(n59), .Z(\ab[13][9] ) );
  NR2 U1100 ( .A(n21), .B(n59), .Z(\ab[13][8] ) );
  NR2 U1101 ( .A(n20), .B(n59), .Z(\ab[13][7] ) );
  NR2 U1102 ( .A(n19), .B(n59), .Z(\ab[13][6] ) );
  NR2 U1103 ( .A(n18), .B(n59), .Z(\ab[13][5] ) );
  NR2 U1104 ( .A(n17), .B(n59), .Z(\ab[13][4] ) );
  NR2 U1105 ( .A(n16), .B(n59), .Z(\ab[13][3] ) );
  NR2 U1106 ( .A(n15), .B(n59), .Z(\ab[13][2] ) );
  NR2 U1107 ( .A(n5), .B(n59), .Z(\ab[13][21] ) );
  NR2 U1108 ( .A(n6), .B(n59), .Z(\ab[13][20] ) );
  NR2 U1109 ( .A(n14), .B(n59), .Z(\ab[13][1] ) );
  NR2 U1110 ( .A(n7), .B(n59), .Z(\ab[13][19] ) );
  NR2 U1111 ( .A(n8), .B(n59), .Z(\ab[13][18] ) );
  NR2 U1112 ( .A(n9), .B(n59), .Z(\ab[13][17] ) );
  NR2 U1113 ( .A(n10), .B(n59), .Z(\ab[13][16] ) );
  NR2 U1114 ( .A(n11), .B(n59), .Z(\ab[13][15] ) );
  NR2 U1115 ( .A(n4), .B(n59), .Z(\ab[13][14] ) );
  NR2 U1116 ( .A(n12), .B(n59), .Z(\ab[13][13] ) );
  NR2 U1117 ( .A(n25), .B(n59), .Z(\ab[13][12] ) );
  NR2 U1118 ( .A(n24), .B(n59), .Z(\ab[13][11] ) );
  NR2 U1119 ( .A(n23), .B(n59), .Z(\ab[13][10] ) );
  NR2 U1120 ( .A(n13), .B(n59), .Z(\ab[13][0] ) );
  NR2 U1121 ( .A(n22), .B(n60), .Z(\ab[12][9] ) );
  NR2 U1122 ( .A(n21), .B(n60), .Z(\ab[12][8] ) );
  NR2 U1123 ( .A(n20), .B(n60), .Z(\ab[12][7] ) );
  NR2 U1124 ( .A(n19), .B(n60), .Z(\ab[12][6] ) );
  NR2 U1125 ( .A(n18), .B(n60), .Z(\ab[12][5] ) );
  NR2 U1126 ( .A(n17), .B(n60), .Z(\ab[12][4] ) );
  NR2 U1127 ( .A(n16), .B(n60), .Z(\ab[12][3] ) );
  NR2 U1128 ( .A(n15), .B(n60), .Z(\ab[12][2] ) );
  NR2 U1129 ( .A(n5), .B(n60), .Z(\ab[12][21] ) );
  NR2 U1130 ( .A(n6), .B(n60), .Z(\ab[12][20] ) );
  NR2 U1131 ( .A(n14), .B(n60), .Z(\ab[12][1] ) );
  NR2 U1132 ( .A(n7), .B(n60), .Z(\ab[12][19] ) );
  NR2 U1133 ( .A(n8), .B(n60), .Z(\ab[12][18] ) );
  NR2 U1134 ( .A(n9), .B(n60), .Z(\ab[12][17] ) );
  NR2 U1135 ( .A(n10), .B(n60), .Z(\ab[12][16] ) );
  NR2 U1136 ( .A(n11), .B(n60), .Z(\ab[12][15] ) );
  NR2 U1137 ( .A(n4), .B(n60), .Z(\ab[12][14] ) );
  NR2 U1138 ( .A(n12), .B(n60), .Z(\ab[12][13] ) );
  NR2 U1139 ( .A(n25), .B(n60), .Z(\ab[12][12] ) );
  NR2 U1140 ( .A(n24), .B(n60), .Z(\ab[12][11] ) );
  NR2 U1141 ( .A(n23), .B(n60), .Z(\ab[12][10] ) );
  NR2 U1142 ( .A(n13), .B(n60), .Z(\ab[12][0] ) );
  NR2 U1143 ( .A(n22), .B(n61), .Z(\ab[11][9] ) );
  NR2 U1144 ( .A(n21), .B(n61), .Z(\ab[11][8] ) );
  NR2 U1145 ( .A(n20), .B(n61), .Z(\ab[11][7] ) );
  NR2 U1146 ( .A(n19), .B(n61), .Z(\ab[11][6] ) );
  NR2 U1147 ( .A(n18), .B(n61), .Z(\ab[11][5] ) );
  NR2 U1148 ( .A(n17), .B(n61), .Z(\ab[11][4] ) );
  NR2 U1149 ( .A(n16), .B(n61), .Z(\ab[11][3] ) );
  NR2 U1150 ( .A(n15), .B(n61), .Z(\ab[11][2] ) );
  NR2 U1151 ( .A(n5), .B(n61), .Z(\ab[11][21] ) );
  NR2 U1152 ( .A(n6), .B(n61), .Z(\ab[11][20] ) );
  NR2 U1153 ( .A(n14), .B(n61), .Z(\ab[11][1] ) );
  NR2 U1154 ( .A(n7), .B(n61), .Z(\ab[11][19] ) );
  NR2 U1155 ( .A(n8), .B(n61), .Z(\ab[11][18] ) );
  NR2 U1156 ( .A(n9), .B(n61), .Z(\ab[11][17] ) );
  NR2 U1157 ( .A(n10), .B(n61), .Z(\ab[11][16] ) );
  NR2 U1158 ( .A(n11), .B(n61), .Z(\ab[11][15] ) );
  NR2 U1159 ( .A(n4), .B(n61), .Z(\ab[11][14] ) );
  NR2 U1160 ( .A(n12), .B(n61), .Z(\ab[11][13] ) );
  NR2 U1161 ( .A(n25), .B(n61), .Z(\ab[11][12] ) );
  NR2 U1162 ( .A(n24), .B(n61), .Z(\ab[11][11] ) );
  NR2 U1163 ( .A(n23), .B(n61), .Z(\ab[11][10] ) );
  NR2 U1164 ( .A(n13), .B(n61), .Z(\ab[11][0] ) );
  NR2 U1165 ( .A(n22), .B(n62), .Z(\ab[10][9] ) );
  NR2 U1166 ( .A(n21), .B(n62), .Z(\ab[10][8] ) );
  NR2 U1167 ( .A(n20), .B(n62), .Z(\ab[10][7] ) );
  NR2 U1168 ( .A(n19), .B(n62), .Z(\ab[10][6] ) );
  NR2 U1169 ( .A(n18), .B(n62), .Z(\ab[10][5] ) );
  NR2 U1170 ( .A(n17), .B(n62), .Z(\ab[10][4] ) );
  NR2 U1171 ( .A(n16), .B(n62), .Z(\ab[10][3] ) );
  NR2 U1172 ( .A(n15), .B(n62), .Z(\ab[10][2] ) );
  NR2 U1173 ( .A(n5), .B(n62), .Z(\ab[10][21] ) );
  NR2 U1174 ( .A(n6), .B(n62), .Z(\ab[10][20] ) );
  NR2 U1175 ( .A(n14), .B(n62), .Z(\ab[10][1] ) );
  NR2 U1176 ( .A(n7), .B(n62), .Z(\ab[10][19] ) );
  NR2 U1177 ( .A(n8), .B(n62), .Z(\ab[10][18] ) );
  NR2 U1178 ( .A(n9), .B(n62), .Z(\ab[10][17] ) );
  NR2 U1179 ( .A(n10), .B(n62), .Z(\ab[10][16] ) );
  NR2 U1180 ( .A(n11), .B(n62), .Z(\ab[10][15] ) );
  NR2 U1181 ( .A(n4), .B(n62), .Z(\ab[10][14] ) );
  NR2 U1182 ( .A(n12), .B(n62), .Z(\ab[10][13] ) );
  NR2 U1183 ( .A(n25), .B(n62), .Z(\ab[10][12] ) );
  NR2 U1184 ( .A(n24), .B(n62), .Z(\ab[10][11] ) );
  NR2 U1185 ( .A(n23), .B(n62), .Z(\ab[10][10] ) );
  NR2 U1186 ( .A(n13), .B(n62), .Z(\ab[10][0] ) );
  NR2 U1187 ( .A(n22), .B(n72), .Z(\ab[0][9] ) );
  NR2 U1188 ( .A(n21), .B(n72), .Z(\ab[0][8] ) );
  NR2 U1189 ( .A(n20), .B(n72), .Z(\ab[0][7] ) );
  NR2 U1190 ( .A(n19), .B(n72), .Z(\ab[0][6] ) );
  NR2 U1191 ( .A(n18), .B(n72), .Z(\ab[0][5] ) );
  NR2 U1192 ( .A(n17), .B(n72), .Z(\ab[0][4] ) );
  NR2 U1193 ( .A(n16), .B(n72), .Z(\ab[0][3] ) );
  NR2 U1194 ( .A(n15), .B(n72), .Z(\ab[0][2] ) );
  NR2 U1195 ( .A(n5), .B(n72), .Z(\ab[0][21] ) );
  NR2 U1196 ( .A(n6), .B(n72), .Z(\ab[0][20] ) );
  NR2 U1197 ( .A(n7), .B(n72), .Z(\ab[0][19] ) );
  NR2 U1198 ( .A(n8), .B(n72), .Z(\ab[0][18] ) );
  NR2 U1199 ( .A(n9), .B(n72), .Z(\ab[0][17] ) );
  NR2 U1200 ( .A(n10), .B(n72), .Z(\ab[0][16] ) );
  NR2 U1201 ( .A(n11), .B(n72), .Z(\ab[0][15] ) );
  NR2 U1202 ( .A(n4), .B(n72), .Z(\ab[0][14] ) );
  NR2 U1203 ( .A(n12), .B(n72), .Z(\ab[0][13] ) );
  NR2 U1204 ( .A(n25), .B(n72), .Z(\ab[0][12] ) );
  NR2 U1205 ( .A(n24), .B(n72), .Z(\ab[0][11] ) );
  NR2 U1206 ( .A(n23), .B(n72), .Z(\ab[0][10] ) );
  AN3 U1207 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U1208 ( .A(n71), .B(n14), .Z(\ab[1][1] ) );
endmodule


module Poly_Logarithm ( clock, reset, input_log, output_log );
  input [47:0] input_log;
  output [30:0] output_log;
  input clock, reset;
  wire   N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N136, N137, N138, N139, N140, N141, N142, n216, n217, n218, n220,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235;
  wire   [47:0] input_log2;
  wire   [67:38] num2;
  wire   [26:1] num3;
  wire   [67:61] num2_1;
  wire   [26:24] num3_1;
  wire   [23:0] Fraction_bit;
  wire   [6:0] Integer_bit;
  wire   [22:0] Log_P;
  wire   [29:0] Log;
  tri   clock;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39;
  assign output_log[0] = 1'b0;

  Poly_Logarithm_DW01_sub_1 sub_0_root_add_364 ( .A({1'b0, N96, N95, N94, N93, 
        N92, N91, N90, N89, N88, N87, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, num2[60:38]}), .CI(
        1'b0), .DIFF({N121, N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, 
        N100, N99, N98}) );
  Poly_Logarithm_DW02_mult_0 mult_357 ( .A(input_log2), .B({n216, n217, n218, 
        n226, n227, n228, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, 
        N25, N26, N27, N28, N29, N30}), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}) );
  FDS2L \num2_1_reg[67]  ( .CR(1'b1), .D(num2[67]), .LD(n2235), .CP(clock), 
        .QN(n2234) );
  FDS2L \Fraction_bit_reg[23]  ( .CR(1'b1), .D(N121), .LD(n2235), .CP(clock), 
        .Q(n229) );
  FDS2L \num3_reg[23]  ( .CR(1'b1), .D(N64), .LD(n2235), .CP(clock), .Q(N96)
         );
  FDS2L \num3_reg[22]  ( .CR(1'b1), .D(N65), .LD(n2235), .CP(clock), .Q(N95)
         );
  FDS2L \num3_reg[21]  ( .CR(1'b1), .D(N66), .LD(n2235), .CP(clock), .Q(N94)
         );
  FDS2L \num3_reg[20]  ( .CR(1'b1), .D(N67), .LD(n2235), .CP(clock), .Q(N93)
         );
  FDS2L \num3_reg[19]  ( .CR(1'b1), .D(N68), .LD(n2235), .CP(clock), .Q(N92)
         );
  FDS2L \num3_reg[18]  ( .CR(1'b1), .D(N69), .LD(n2235), .CP(clock), .Q(N91)
         );
  FDS2L \num3_reg[17]  ( .CR(1'b1), .D(N70), .LD(n2235), .CP(clock), .Q(N90)
         );
  FDS2L \num3_reg[16]  ( .CR(1'b1), .D(N71), .LD(n2235), .CP(clock), .Q(N89)
         );
  FDS2L \num3_reg[15]  ( .CR(1'b1), .D(N72), .LD(n2235), .CP(clock), .Q(N88)
         );
  FDS2L \num3_reg[14]  ( .CR(1'b1), .D(N73), .LD(n2235), .CP(clock), .Q(N87)
         );
  FDS2L \num2_1_reg[65]  ( .CR(1'b1), .D(num2[65]), .LD(n2235), .CP(clock), 
        .Q(num2_1[65]), .QN(n230) );
  FDS2L \num2_1_reg[63]  ( .CR(1'b1), .D(num2[63]), .LD(n2235), .CP(clock), 
        .Q(num2_1[63]) );
  FDS2L \num2_1_reg[62]  ( .CR(1'b1), .D(num2[62]), .LD(n2235), .CP(clock), 
        .Q(num2_1[62]) );
  FDS2L \num2_1_reg[61]  ( .CR(1'b1), .D(num2[61]), .LD(n2235), .CP(clock), 
        .Q(num2_1[61]) );
  FDS2L \input_log2_reg[39]  ( .CR(1'b1), .D(input_log[39]), .LD(n2235), .CP(
        clock), .Q(input_log2[39]) );
  FDS2L \input_log2_reg[38]  ( .CR(1'b1), .D(input_log[38]), .LD(n2235), .CP(
        clock), .Q(input_log2[38]) );
  FDS2L \input_log2_reg[37]  ( .CR(1'b1), .D(input_log[37]), .LD(n2235), .CP(
        clock), .Q(input_log2[37]) );
  FDS2L \input_log2_reg[36]  ( .CR(1'b1), .D(input_log[36]), .LD(n2235), .CP(
        clock), .Q(input_log2[36]) );
  FDS2L \input_log2_reg[35]  ( .CR(1'b1), .D(input_log[35]), .LD(n2235), .CP(
        clock), .Q(input_log2[35]) );
  FDS2L \input_log2_reg[34]  ( .CR(1'b1), .D(input_log[34]), .LD(n2235), .CP(
        clock), .Q(input_log2[34]) );
  FDS2L \input_log2_reg[33]  ( .CR(1'b1), .D(input_log[33]), .LD(n2235), .CP(
        clock), .Q(input_log2[33]) );
  FDS2L \input_log2_reg[32]  ( .CR(1'b1), .D(input_log[32]), .LD(n2235), .CP(
        clock), .Q(input_log2[32]) );
  FDS2L \input_log2_reg[31]  ( .CR(1'b1), .D(input_log[31]), .LD(n2235), .CP(
        clock), .Q(input_log2[31]) );
  FDS2L \input_log2_reg[30]  ( .CR(1'b1), .D(input_log[30]), .LD(n2235), .CP(
        clock), .Q(input_log2[30]) );
  FDS2L \input_log2_reg[29]  ( .CR(1'b1), .D(input_log[29]), .LD(n2235), .CP(
        clock), .Q(input_log2[29]) );
  FDS2L \input_log2_reg[28]  ( .CR(1'b1), .D(input_log[28]), .LD(n2235), .CP(
        clock), .Q(input_log2[28]) );
  FDS2L \input_log2_reg[27]  ( .CR(1'b1), .D(input_log[27]), .LD(n2235), .CP(
        clock), .Q(input_log2[27]) );
  FDS2L \input_log2_reg[26]  ( .CR(1'b1), .D(input_log[26]), .LD(n2235), .CP(
        clock), .Q(input_log2[26]) );
  FDS2L \input_log2_reg[25]  ( .CR(1'b1), .D(input_log[25]), .LD(n2235), .CP(
        clock), .Q(input_log2[25]) );
  FDS2L \input_log2_reg[24]  ( .CR(1'b1), .D(input_log[24]), .LD(n2235), .CP(
        clock), .Q(input_log2[24]) );
  FDS2L \input_log2_reg[23]  ( .CR(1'b1), .D(input_log[23]), .LD(n2235), .CP(
        clock), .Q(input_log2[23]) );
  FDS2L \input_log2_reg[22]  ( .CR(1'b1), .D(input_log[22]), .LD(n2235), .CP(
        clock), .Q(input_log2[22]) );
  FDS2L \input_log2_reg[21]  ( .CR(1'b1), .D(input_log[21]), .LD(n2235), .CP(
        clock), .Q(input_log2[21]) );
  FDS2L \input_log2_reg[20]  ( .CR(1'b1), .D(input_log[20]), .LD(n2235), .CP(
        clock), .Q(input_log2[20]) );
  FDS2L \input_log2_reg[19]  ( .CR(1'b1), .D(input_log[19]), .LD(n2235), .CP(
        clock), .Q(input_log2[19]) );
  FDS2L \input_log2_reg[18]  ( .CR(1'b1), .D(input_log[18]), .LD(n2235), .CP(
        clock), .Q(input_log2[18]) );
  FDS2L \input_log2_reg[17]  ( .CR(1'b1), .D(input_log[17]), .LD(n2235), .CP(
        clock), .Q(input_log2[17]) );
  FDS2L \input_log2_reg[16]  ( .CR(1'b1), .D(input_log[16]), .LD(n2235), .CP(
        clock), .Q(input_log2[16]) );
  FDS2L \input_log2_reg[15]  ( .CR(1'b1), .D(input_log[15]), .LD(n2235), .CP(
        clock), .Q(input_log2[15]) );
  FDS2L \input_log2_reg[14]  ( .CR(1'b1), .D(input_log[14]), .LD(n2235), .CP(
        clock), .Q(input_log2[14]) );
  FDS2L \input_log2_reg[13]  ( .CR(1'b1), .D(input_log[13]), .LD(n2235), .CP(
        clock), .Q(input_log2[13]) );
  FDS2L \input_log2_reg[12]  ( .CR(1'b1), .D(input_log[12]), .LD(n2235), .CP(
        clock), .Q(input_log2[12]) );
  FDS2L \input_log2_reg[11]  ( .CR(1'b1), .D(input_log[11]), .LD(n2235), .CP(
        clock), .Q(input_log2[11]) );
  FDS2L \input_log2_reg[10]  ( .CR(1'b1), .D(input_log[10]), .LD(n2235), .CP(
        clock), .Q(input_log2[10]) );
  FDS2L \input_log2_reg[9]  ( .CR(1'b1), .D(input_log[9]), .LD(n2235), .CP(
        clock), .Q(input_log2[9]) );
  FDS2L \input_log2_reg[8]  ( .CR(1'b1), .D(input_log[8]), .LD(n2235), .CP(
        clock), .Q(input_log2[8]) );
  FDS2L \input_log2_reg[7]  ( .CR(1'b1), .D(input_log[7]), .LD(n2235), .CP(
        clock), .Q(input_log2[7]) );
  FDS2L \input_log2_reg[6]  ( .CR(1'b1), .D(input_log[6]), .LD(n2235), .CP(
        clock), .Q(input_log2[6]) );
  FDS2L \input_log2_reg[5]  ( .CR(1'b1), .D(input_log[5]), .LD(n2235), .CP(
        clock), .Q(input_log2[5]) );
  FDS2L \input_log2_reg[4]  ( .CR(1'b1), .D(input_log[4]), .LD(n2235), .CP(
        clock), .Q(input_log2[4]) );
  FDS2L \input_log2_reg[3]  ( .CR(1'b1), .D(input_log[3]), .LD(n2235), .CP(
        clock), .Q(input_log2[3]) );
  FDS2L \input_log2_reg[2]  ( .CR(1'b1), .D(input_log[2]), .LD(n2235), .CP(
        clock), .Q(input_log2[2]) );
  FDS2L \input_log2_reg[1]  ( .CR(1'b1), .D(input_log[1]), .LD(n2235), .CP(
        clock), .Q(input_log2[1]) );
  FDS2L \num2_reg[60]  ( .CR(1'b1), .D(N53), .LD(n2235), .CP(clock), .Q(
        num2[60]) );
  FDS2L \num2_reg[59]  ( .CR(1'b1), .D(N52), .LD(n2235), .CP(clock), .Q(
        num2[59]) );
  FDS2L \num2_reg[58]  ( .CR(1'b1), .D(N51), .LD(n2235), .CP(clock), .Q(
        num2[58]) );
  FDS2L \num2_reg[57]  ( .CR(1'b1), .D(N50), .LD(n2235), .CP(clock), .Q(
        num2[57]) );
  FDS2L \num2_reg[56]  ( .CR(1'b1), .D(N49), .LD(n2235), .CP(clock), .Q(
        num2[56]) );
  FDS2L \num2_reg[55]  ( .CR(1'b1), .D(N48), .LD(n2235), .CP(clock), .Q(
        num2[55]) );
  FDS2L \num2_reg[54]  ( .CR(1'b1), .D(N47), .LD(n2235), .CP(clock), .Q(
        num2[54]) );
  FDS2L \num2_reg[53]  ( .CR(1'b1), .D(N46), .LD(n2235), .CP(clock), .Q(
        num2[53]) );
  FDS2L \num2_reg[52]  ( .CR(1'b1), .D(N45), .LD(n2235), .CP(clock), .Q(
        num2[52]) );
  FDS2L \num2_reg[51]  ( .CR(1'b1), .D(N44), .LD(n2235), .CP(clock), .Q(
        num2[51]) );
  FDS2L \num2_reg[50]  ( .CR(1'b1), .D(N43), .LD(n2235), .CP(clock), .Q(
        num2[50]) );
  FDS2L \num2_reg[49]  ( .CR(1'b1), .D(N42), .LD(n2235), .CP(clock), .Q(
        num2[49]) );
  FDS2L \num2_reg[48]  ( .CR(1'b1), .D(N41), .LD(n2235), .CP(clock), .Q(
        num2[48]) );
  FDS2L \num2_reg[47]  ( .CR(1'b1), .D(N40), .LD(n2235), .CP(clock), .Q(
        num2[47]) );
  FDS2L \num2_reg[46]  ( .CR(1'b1), .D(N39), .LD(n2235), .CP(clock), .Q(
        num2[46]) );
  FDS2L \num2_reg[45]  ( .CR(1'b1), .D(N38), .LD(n2235), .CP(clock), .Q(
        num2[45]) );
  FDS2L \num2_reg[44]  ( .CR(1'b1), .D(N37), .LD(n2235), .CP(clock), .Q(
        num2[44]) );
  FDS2L \num2_reg[43]  ( .CR(1'b1), .D(N36), .LD(n2235), .CP(clock), .Q(
        num2[43]) );
  FDS2L \num2_reg[42]  ( .CR(1'b1), .D(N35), .LD(n2235), .CP(clock), .Q(
        num2[42]) );
  FDS2L \num2_reg[41]  ( .CR(1'b1), .D(N34), .LD(n2235), .CP(clock), .Q(
        num2[41]) );
  FDS2L \num2_reg[40]  ( .CR(1'b1), .D(N33), .LD(n2235), .CP(clock), .Q(
        num2[40]) );
  FDS2L \num2_reg[39]  ( .CR(1'b1), .D(N32), .LD(n2235), .CP(clock), .Q(
        num2[39]) );
  FDS2L \num2_1_reg[66]  ( .CR(1'b1), .D(num2[66]), .LD(n2235), .CP(clock), 
        .Q(num2_1[66]) );
  FDS2L \num2_1_reg[64]  ( .CR(1'b1), .D(num2[64]), .LD(n2235), .CP(clock), 
        .Q(num2_1[64]) );
  FDS2L \num3_1_reg[26]  ( .CR(1'b1), .D(num3[26]), .LD(n2235), .CP(clock), 
        .Q(num3_1[26]) );
  FDS2L \num3_1_reg[25]  ( .CR(1'b1), .D(num3[25]), .LD(n2235), .CP(clock), 
        .Q(num3_1[25]) );
  FDS2L \output_log_reg[24]  ( .CR(1'b1), .D(Log[23]), .LD(n2235), .CP(clock), 
        .Q(output_log[24]) );
  FDS2L \output_log_reg[23]  ( .CR(1'b1), .D(Log[22]), .LD(n2235), .CP(clock), 
        .Q(output_log[23]) );
  FDS2L \output_log_reg[22]  ( .CR(1'b1), .D(Log[21]), .LD(n2235), .CP(clock), 
        .Q(output_log[22]) );
  FDS2L \output_log_reg[21]  ( .CR(1'b1), .D(Log[20]), .LD(n2235), .CP(clock), 
        .Q(output_log[21]) );
  FDS2L \output_log_reg[20]  ( .CR(1'b1), .D(Log[19]), .LD(n2235), .CP(clock), 
        .Q(output_log[20]) );
  FDS2L \output_log_reg[19]  ( .CR(1'b1), .D(Log[18]), .LD(n2235), .CP(clock), 
        .Q(output_log[19]) );
  FDS2L \output_log_reg[18]  ( .CR(1'b1), .D(Log[17]), .LD(n2235), .CP(clock), 
        .Q(output_log[18]) );
  FDS2L \output_log_reg[17]  ( .CR(1'b1), .D(Log[16]), .LD(n2235), .CP(clock), 
        .Q(output_log[17]) );
  FDS2L \output_log_reg[16]  ( .CR(1'b1), .D(Log[15]), .LD(n2235), .CP(clock), 
        .Q(output_log[16]) );
  FDS2L \output_log_reg[15]  ( .CR(1'b1), .D(Log[14]), .LD(n2235), .CP(clock), 
        .Q(output_log[15]) );
  FDS2L \output_log_reg[14]  ( .CR(1'b1), .D(Log[13]), .LD(n2235), .CP(clock), 
        .Q(output_log[14]) );
  FDS2L \output_log_reg[13]  ( .CR(1'b1), .D(Log[12]), .LD(n2235), .CP(clock), 
        .Q(output_log[13]) );
  FDS2L \output_log_reg[12]  ( .CR(1'b1), .D(Log[11]), .LD(n2235), .CP(clock), 
        .Q(output_log[12]) );
  FDS2L \output_log_reg[11]  ( .CR(1'b1), .D(Log[10]), .LD(n2235), .CP(clock), 
        .Q(output_log[11]) );
  FDS2L \output_log_reg[10]  ( .CR(1'b1), .D(Log[9]), .LD(n2235), .CP(clock), 
        .Q(output_log[10]) );
  FDS2L \output_log_reg[9]  ( .CR(1'b1), .D(Log[8]), .LD(n2235), .CP(clock), 
        .Q(output_log[9]) );
  FDS2L \output_log_reg[8]  ( .CR(1'b1), .D(Log[7]), .LD(n2235), .CP(clock), 
        .Q(output_log[8]) );
  FDS2L \output_log_reg[7]  ( .CR(1'b1), .D(Log[6]), .LD(n2235), .CP(clock), 
        .Q(output_log[7]) );
  FDS2L \output_log_reg[6]  ( .CR(1'b1), .D(Log[5]), .LD(n2235), .CP(clock), 
        .Q(output_log[6]) );
  FDS2L \output_log_reg[5]  ( .CR(1'b1), .D(Log[4]), .LD(n2235), .CP(clock), 
        .Q(output_log[5]) );
  FDS2L \output_log_reg[4]  ( .CR(1'b1), .D(Log[3]), .LD(n2235), .CP(clock), 
        .Q(output_log[4]) );
  FDS2L \output_log_reg[3]  ( .CR(1'b1), .D(Log[2]), .LD(n2235), .CP(clock), 
        .Q(output_log[3]) );
  FDS2L \output_log_reg[2]  ( .CR(1'b1), .D(Log[1]), .LD(n2235), .CP(clock), 
        .Q(output_log[2]) );
  FDS2L \output_log_reg[1]  ( .CR(1'b1), .D(Log[0]), .LD(n2235), .CP(clock), 
        .Q(output_log[1]) );
  FDS2L \input_log2_reg[0]  ( .CR(1'b1), .D(input_log[0]), .LD(n2235), .CP(
        clock), .Q(input_log2[0]) );
  FDS2L \num2_reg[38]  ( .CR(1'b1), .D(N31), .LD(n2235), .CP(clock), .Q(
        num2[38]) );
  FDS2L \num3_1_reg[24]  ( .CR(1'b1), .D(num3[24]), .LD(n2235), .CP(clock), 
        .Q(num3_1[24]) );
  FDS2L \output_log_reg[30]  ( .CR(1'b1), .D(Log[29]), .LD(n2235), .CP(clock), 
        .Q(output_log[30]) );
  FDS2L \input_log2_reg[46]  ( .CR(1'b1), .D(input_log[46]), .LD(n2235), .CP(
        clock), .Q(input_log2[46]), .QN(n222) );
  FDS2L \output_log_reg[28]  ( .CR(1'b1), .D(Log[27]), .LD(n2235), .CP(clock), 
        .Q(output_log[28]) );
  FDS2L \input_log2_reg[47]  ( .CR(1'b1), .D(input_log[47]), .LD(n2235), .CP(
        clock), .Q(input_log2[47]), .QN(n220) );
  FDS2L \output_log_reg[29]  ( .CR(1'b1), .D(Log[28]), .LD(n2235), .CP(clock), 
        .Q(output_log[29]) );
  FDS2L \output_log_reg[26]  ( .CR(1'b1), .D(Log[25]), .LD(n2235), .CP(clock), 
        .Q(output_log[26]) );
  FDS2L \output_log_reg[25]  ( .CR(1'b1), .D(Log[24]), .LD(n2235), .CP(clock), 
        .Q(output_log[25]) );
  FDS2L \input_log2_reg[45]  ( .CR(1'b1), .D(input_log[45]), .LD(n2235), .CP(
        clock), .Q(input_log2[45]), .QN(n278) );
  FDS2L \output_log_reg[27]  ( .CR(1'b1), .D(Log[26]), .LD(n2235), .CP(clock), 
        .Q(output_log[27]) );
  FDS2L \input_log2_reg[43]  ( .CR(1'b1), .D(input_log[43]), .LD(n2235), .CP(
        clock), .Q(input_log2[43]), .QN(n277) );
  FDS2L \input_log2_reg[44]  ( .CR(1'b1), .D(input_log[44]), .LD(n2235), .CP(
        clock), .Q(input_log2[44]), .QN(n279) );
  FDS2L \input_log2_reg[40]  ( .CR(1'b1), .D(input_log[40]), .LD(n2235), .CP(
        clock), .Q(input_log2[40]), .QN(n225) );
  FDS2L \input_log2_reg[41]  ( .CR(1'b1), .D(input_log[41]), .LD(n2235), .CP(
        clock), .Q(input_log2[41]), .QN(n224) );
  FDS2L \input_log2_reg[42]  ( .CR(1'b1), .D(input_log[42]), .LD(n2235), .CP(
        clock), .Q(input_log2[42]), .QN(n223) );
  FDS2L \num2_reg[67]  ( .CR(1'b1), .D(N60), .LD(n2235), .CP(clock), .Q(
        num2[67]) );
  FDS2L \num2_reg[66]  ( .CR(1'b1), .D(N59), .LD(n2235), .CP(clock), .Q(
        num2[66]) );
  FDS2L \num2_reg[65]  ( .CR(1'b1), .D(N58), .LD(n2235), .CP(clock), .Q(
        num2[65]) );
  FDS2L \num2_reg[64]  ( .CR(1'b1), .D(N57), .LD(n2235), .CP(clock), .Q(
        num2[64]) );
  FDS2L \num2_reg[63]  ( .CR(1'b1), .D(N56), .LD(n2235), .CP(clock), .Q(
        num2[63]) );
  FDS2L \num2_reg[62]  ( .CR(1'b1), .D(N55), .LD(n2235), .CP(clock), .Q(
        num2[62]) );
  FDS2L \num2_reg[61]  ( .CR(1'b1), .D(N54), .LD(n2235), .CP(clock), .Q(
        num2[61]) );
  FDS2L \num3_reg[26]  ( .CR(1'b1), .D(n239), .LD(n2235), .CP(clock), .Q(
        num3[26]) );
  FDS2L \num3_reg[25]  ( .CR(1'b1), .D(N62), .LD(n2235), .CP(clock), .Q(
        num3[25]) );
  FDS2L \num3_reg[24]  ( .CR(1'b1), .D(N63), .LD(n2235), .CP(clock), .Q(
        num3[24]) );
  FDS2L \Fraction_bit_reg[22]  ( .CR(1'b1), .D(N120), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[22]) );
  FDS2L \Fraction_bit_reg[21]  ( .CR(1'b1), .D(N119), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[21]) );
  FDS2L \Fraction_bit_reg[20]  ( .CR(1'b1), .D(N118), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[20]) );
  FDS2L \Fraction_bit_reg[19]  ( .CR(1'b1), .D(N117), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[19]) );
  FDS2L \Fraction_bit_reg[18]  ( .CR(1'b1), .D(N116), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[18]) );
  FDS2L \Fraction_bit_reg[17]  ( .CR(1'b1), .D(N115), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[17]) );
  FDS2L \Fraction_bit_reg[16]  ( .CR(1'b1), .D(N114), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[16]) );
  FDS2L \Fraction_bit_reg[15]  ( .CR(1'b1), .D(N113), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[15]) );
  FDS2L \Fraction_bit_reg[14]  ( .CR(1'b1), .D(N112), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[14]) );
  FDS2L \Fraction_bit_reg[13]  ( .CR(1'b1), .D(N111), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[13]) );
  FDS2L \Fraction_bit_reg[12]  ( .CR(1'b1), .D(N110), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[12]) );
  FDS2L \Fraction_bit_reg[11]  ( .CR(1'b1), .D(N109), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[11]) );
  FDS2L \Fraction_bit_reg[10]  ( .CR(1'b1), .D(N108), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[10]) );
  FDS2L \Fraction_bit_reg[9]  ( .CR(1'b1), .D(N107), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[9]) );
  FDS2L \Fraction_bit_reg[8]  ( .CR(1'b1), .D(N106), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[8]) );
  FDS2L \Fraction_bit_reg[7]  ( .CR(1'b1), .D(N105), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[7]) );
  FDS2L \Fraction_bit_reg[6]  ( .CR(1'b1), .D(N104), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[6]) );
  FDS2L \Fraction_bit_reg[5]  ( .CR(1'b1), .D(N103), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[5]) );
  FDS2L \Fraction_bit_reg[4]  ( .CR(1'b1), .D(N102), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[4]) );
  FDS2L \Fraction_bit_reg[3]  ( .CR(1'b1), .D(N101), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[3]) );
  FDS2L \Fraction_bit_reg[2]  ( .CR(1'b1), .D(N100), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[2]) );
  FDS2L \Fraction_bit_reg[1]  ( .CR(1'b1), .D(N99), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[1]) );
  FDS2L \Fraction_bit_reg[0]  ( .CR(1'b1), .D(N98), .LD(n2235), .CP(clock), 
        .Q(Fraction_bit[0]) );
  FDS2L \Integer_bit_reg[6]  ( .CR(1'b1), .D(N142), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[6]) );
  FDS2L \Integer_bit_reg[5]  ( .CR(1'b1), .D(N141), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[5]) );
  FDS2L \Integer_bit_reg[4]  ( .CR(1'b1), .D(N140), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[4]) );
  FDS2L \Integer_bit_reg[3]  ( .CR(1'b1), .D(N139), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[3]) );
  FDS2L \Integer_bit_reg[2]  ( .CR(1'b1), .D(N138), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[2]) );
  FDS2L \Integer_bit_reg[1]  ( .CR(1'b1), .D(N137), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[1]) );
  FDS2L \Integer_bit_reg[0]  ( .CR(1'b1), .D(N136), .LD(n2235), .CP(clock), 
        .Q(Integer_bit[0]) );
  FDS2L \Log_P_reg[22]  ( .CR(1'b1), .D(Fraction_bit[22]), .LD(n2235), .CP(
        clock), .Q(Log_P[22]) );
  FDS2L \Log_P_reg[21]  ( .CR(1'b1), .D(Fraction_bit[21]), .LD(n2235), .CP(
        clock), .Q(Log_P[21]) );
  FDS2L \Log_P_reg[20]  ( .CR(1'b1), .D(Fraction_bit[20]), .LD(n2235), .CP(
        clock), .Q(Log_P[20]) );
  FDS2L \Log_P_reg[19]  ( .CR(1'b1), .D(Fraction_bit[19]), .LD(n2235), .CP(
        clock), .Q(Log_P[19]) );
  FDS2L \Log_P_reg[18]  ( .CR(1'b1), .D(Fraction_bit[18]), .LD(n2235), .CP(
        clock), .Q(Log_P[18]) );
  FDS2L \Log_P_reg[17]  ( .CR(1'b1), .D(Fraction_bit[17]), .LD(n2235), .CP(
        clock), .Q(Log_P[17]) );
  FDS2L \Log_P_reg[16]  ( .CR(1'b1), .D(Fraction_bit[16]), .LD(n2235), .CP(
        clock), .Q(Log_P[16]) );
  FDS2L \Log_P_reg[15]  ( .CR(1'b1), .D(Fraction_bit[15]), .LD(n2235), .CP(
        clock), .Q(Log_P[15]) );
  FDS2L \Log_P_reg[14]  ( .CR(1'b1), .D(Fraction_bit[14]), .LD(n2235), .CP(
        clock), .Q(Log_P[14]) );
  FDS2L \Log_P_reg[13]  ( .CR(1'b1), .D(Fraction_bit[13]), .LD(n2235), .CP(
        clock), .Q(Log_P[13]) );
  FDS2L \Log_P_reg[12]  ( .CR(1'b1), .D(Fraction_bit[12]), .LD(n2235), .CP(
        clock), .Q(Log_P[12]) );
  FDS2L \Log_P_reg[11]  ( .CR(1'b1), .D(Fraction_bit[11]), .LD(n2235), .CP(
        clock), .Q(Log_P[11]) );
  FDS2L \Log_P_reg[10]  ( .CR(1'b1), .D(Fraction_bit[10]), .LD(n2235), .CP(
        clock), .Q(Log_P[10]) );
  FDS2L \Log_P_reg[9]  ( .CR(1'b1), .D(Fraction_bit[9]), .LD(n2235), .CP(clock), .Q(Log_P[9]) );
  FDS2L \Log_P_reg[8]  ( .CR(1'b1), .D(Fraction_bit[8]), .LD(n2235), .CP(clock), .Q(Log_P[8]) );
  FDS2L \Log_P_reg[7]  ( .CR(1'b1), .D(Fraction_bit[7]), .LD(n2235), .CP(clock), .Q(Log_P[7]) );
  FDS2L \Log_P_reg[6]  ( .CR(1'b1), .D(Fraction_bit[6]), .LD(n2235), .CP(clock), .Q(Log_P[6]) );
  FDS2L \Log_P_reg[5]  ( .CR(1'b1), .D(Fraction_bit[5]), .LD(n2235), .CP(clock), .Q(Log_P[5]) );
  FDS2L \Log_P_reg[4]  ( .CR(1'b1), .D(Fraction_bit[4]), .LD(n2235), .CP(clock), .Q(Log_P[4]) );
  FDS2L \Log_P_reg[3]  ( .CR(1'b1), .D(Fraction_bit[3]), .LD(n2235), .CP(clock), .Q(Log_P[3]) );
  FDS2L \Log_P_reg[2]  ( .CR(1'b1), .D(Fraction_bit[2]), .LD(n2235), .CP(clock), .Q(Log_P[2]) );
  FDS2L \Log_P_reg[1]  ( .CR(1'b1), .D(Fraction_bit[1]), .LD(n2235), .CP(clock), .Q(Log_P[1]) );
  FDS2L \Log_P_reg[0]  ( .CR(1'b1), .D(Fraction_bit[0]), .LD(n2235), .CP(clock), .Q(Log_P[0]) );
  FDS2L \Log_reg[29]  ( .CR(1'b1), .D(Integer_bit[6]), .LD(n2235), .CP(clock), 
        .Q(Log[29]) );
  FDS2L \Log_reg[28]  ( .CR(1'b1), .D(Integer_bit[5]), .LD(n2235), .CP(clock), 
        .Q(Log[28]) );
  FDS2L \Log_reg[27]  ( .CR(1'b1), .D(Integer_bit[4]), .LD(n2235), .CP(clock), 
        .Q(Log[27]) );
  FDS2L \Log_reg[26]  ( .CR(1'b1), .D(Integer_bit[3]), .LD(n2235), .CP(clock), 
        .Q(Log[26]) );
  FDS2L \Log_reg[25]  ( .CR(1'b1), .D(Integer_bit[2]), .LD(n2235), .CP(clock), 
        .Q(Log[25]) );
  FDS2L \Log_reg[24]  ( .CR(1'b1), .D(Integer_bit[1]), .LD(n2235), .CP(clock), 
        .Q(Log[24]) );
  FDS2L \Log_reg[23]  ( .CR(1'b1), .D(Integer_bit[0]), .LD(n2235), .CP(clock), 
        .Q(Log[23]) );
  FDS2L \Log_reg[22]  ( .CR(1'b1), .D(Log_P[22]), .LD(n2235), .CP(clock), .Q(
        Log[22]) );
  FDS2L \Log_reg[21]  ( .CR(1'b1), .D(Log_P[21]), .LD(n2235), .CP(clock), .Q(
        Log[21]) );
  FDS2L \Log_reg[20]  ( .CR(1'b1), .D(Log_P[20]), .LD(n2235), .CP(clock), .Q(
        Log[20]) );
  FDS2L \Log_reg[19]  ( .CR(1'b1), .D(Log_P[19]), .LD(n2235), .CP(clock), .Q(
        Log[19]) );
  FDS2L \Log_reg[18]  ( .CR(1'b1), .D(Log_P[18]), .LD(n2235), .CP(clock), .Q(
        Log[18]) );
  FDS2L \Log_reg[17]  ( .CR(1'b1), .D(Log_P[17]), .LD(n2235), .CP(clock), .Q(
        Log[17]) );
  FDS2L \Log_reg[16]  ( .CR(1'b1), .D(Log_P[16]), .LD(n2235), .CP(clock), .Q(
        Log[16]) );
  FDS2L \Log_reg[15]  ( .CR(1'b1), .D(Log_P[15]), .LD(n2235), .CP(clock), .Q(
        Log[15]) );
  FDS2L \Log_reg[14]  ( .CR(1'b1), .D(Log_P[14]), .LD(n2235), .CP(clock), .Q(
        Log[14]) );
  FDS2L \Log_reg[13]  ( .CR(1'b1), .D(Log_P[13]), .LD(n2235), .CP(clock), .Q(
        Log[13]) );
  FDS2L \Log_reg[12]  ( .CR(1'b1), .D(Log_P[12]), .LD(n2235), .CP(clock), .Q(
        Log[12]) );
  FDS2L \Log_reg[11]  ( .CR(1'b1), .D(Log_P[11]), .LD(n2235), .CP(clock), .Q(
        Log[11]) );
  FDS2L \Log_reg[10]  ( .CR(1'b1), .D(Log_P[10]), .LD(n2235), .CP(clock), .Q(
        Log[10]) );
  FDS2L \Log_reg[9]  ( .CR(1'b1), .D(Log_P[9]), .LD(n2235), .CP(clock), .Q(
        Log[9]) );
  FDS2L \Log_reg[8]  ( .CR(1'b1), .D(Log_P[8]), .LD(n2235), .CP(clock), .Q(
        Log[8]) );
  FDS2L \Log_reg[7]  ( .CR(1'b1), .D(Log_P[7]), .LD(n2235), .CP(clock), .Q(
        Log[7]) );
  FDS2L \Log_reg[6]  ( .CR(1'b1), .D(Log_P[6]), .LD(n2235), .CP(clock), .Q(
        Log[6]) );
  FDS2L \Log_reg[5]  ( .CR(1'b1), .D(Log_P[5]), .LD(n2235), .CP(clock), .Q(
        Log[5]) );
  FDS2L \Log_reg[4]  ( .CR(1'b1), .D(Log_P[4]), .LD(n2235), .CP(clock), .Q(
        Log[4]) );
  FDS2L \Log_reg[3]  ( .CR(1'b1), .D(Log_P[3]), .LD(n2235), .CP(clock), .Q(
        Log[3]) );
  FDS2L \Log_reg[2]  ( .CR(1'b1), .D(Log_P[2]), .LD(n2235), .CP(clock), .Q(
        Log[2]) );
  FDS2L \Log_reg[1]  ( .CR(1'b1), .D(Log_P[1]), .LD(n2235), .CP(clock), .Q(
        Log[1]) );
  FDS2L \Log_reg[0]  ( .CR(1'b1), .D(Log_P[0]), .LD(n2235), .CP(clock), .Q(
        Log[0]) );
  NR3 U3 ( .A(input_log2[45]), .B(input_log2[43]), .C(n276), .Z(n2070) );
  AN3 U4 ( .A(n220), .B(n222), .C(n238), .Z(n216) );
  AN3 U5 ( .A(n220), .B(n222), .C(n236), .Z(n217) );
  AN3 U6 ( .A(n220), .B(n222), .C(n237), .Z(n218) );
  AN3 U7 ( .A(n220), .B(n222), .C(n560), .Z(n226) );
  AN3 U8 ( .A(n220), .B(n222), .C(n562), .Z(n227) );
  AN3 U9 ( .A(n220), .B(n222), .C(n566), .Z(n228) );
  AN4P U10 ( .A(n312), .B(n278), .C(n279), .D(n277), .Z(n231) );
  AN2P U11 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n232) );
  AN3 U12 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n233) );
  AN3 U13 ( .A(n223), .B(n225), .C(input_log2[41]), .Z(n234) );
  AN2P U14 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n235) );
  AN4P U15 ( .A(n557), .B(n278), .C(n279), .D(n277), .Z(n236) );
  AN4P U16 ( .A(n558), .B(n278), .C(n279), .D(n277), .Z(n237) );
  AN4P U17 ( .A(n556), .B(n278), .C(n279), .D(n277), .Z(n238) );
  AN3 U18 ( .A(n220), .B(n222), .C(n293), .Z(n239) );
  AN2P U19 ( .A(n1752), .B(n1751), .Z(n240) );
  MUX21H U20 ( .A(input_log2[42]), .B(n1111), .S(input_log2[40]), .Z(n241) );
  AN2P U21 ( .A(n1121), .B(n1120), .Z(n242) );
  MUX21H U22 ( .A(n1558), .B(n1557), .S(input_log2[42]), .Z(n243) );
  AN3 U23 ( .A(n1539), .B(n1538), .C(n1537), .Z(n244) );
  AN2P U24 ( .A(n1143), .B(n223), .Z(n245) );
  AN2P U25 ( .A(n1104), .B(n1103), .Z(n246) );
  AN3 U26 ( .A(n1441), .B(n1440), .C(n1439), .Z(n247) );
  MUX21H U27 ( .A(input_log2[41]), .B(input_log2[42]), .S(input_log2[40]), .Z(
        n248) );
  AN2P U28 ( .A(n1127), .B(n1126), .Z(n249) );
  AN3 U29 ( .A(n1130), .B(n1129), .C(n1128), .Z(n250) );
  AN2P U30 ( .A(n1228), .B(n1227), .Z(n251) );
  MUX21H U31 ( .A(n1140), .B(n1139), .S(input_log2[40]), .Z(n252) );
  AN2P U32 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n253) );
  OR3 U33 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n254) );
  AN2P U34 ( .A(n1844), .B(n1843), .Z(n255) );
  AN2P U35 ( .A(n1512), .B(n1511), .Z(n256) );
  AN2P U36 ( .A(n1323), .B(n1322), .Z(n257) );
  AN2P U37 ( .A(n1245), .B(n1244), .Z(n258) );
  AN2P U38 ( .A(n1521), .B(n1520), .Z(n259) );
  AN3 U39 ( .A(input_log2[45]), .B(n1923), .C(n1922), .Z(n260) );
  AN2P U40 ( .A(n1188), .B(n223), .Z(n261) );
  ND3 U41 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .Z(
        n262) );
  OR3 U42 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n263) );
  AN2P U43 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n264) );
  AN2P U44 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n265) );
  AN2P U45 ( .A(n1813), .B(n1812), .Z(n266) );
  AN2P U46 ( .A(n1575), .B(n1574), .Z(n267) );
  AN2P U47 ( .A(n1450), .B(n1449), .Z(n268) );
  MUX21H U48 ( .A(n1502), .B(n1501), .S(input_log2[40]), .Z(n269) );
  MUX21H U49 ( .A(n1329), .B(input_log2[41]), .S(input_log2[42]), .Z(n270) );
  OR2P U50 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n271) );
  AN2P U51 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n272) );
  AN2P U52 ( .A(n1825), .B(n1824), .Z(n273) );
  AN4P U53 ( .A(n2092), .B(n2091), .C(n2090), .D(n2089), .Z(n274) );
  AN4P U54 ( .A(n2102), .B(n2101), .C(n2100), .D(n2099), .Z(n275) );
  ND2 U55 ( .A(n2062), .B(n2061), .Z(n560) );
  ND2 U56 ( .A(n2060), .B(n2059), .Z(n562) );
  AO7 U57 ( .A(n2208), .B(n2007), .C(n2006), .Z(n572) );
  IVP U58 ( .A(n571), .Z(n2208) );
  ND2 U59 ( .A(n278), .B(n277), .Z(n2007) );
  ND2 U60 ( .A(n278), .B(n279), .Z(n2006) );
  ND3 U61 ( .A(n224), .B(n225), .C(n223), .Z(n885) );
  ND3 U62 ( .A(n1367), .B(n1366), .C(n1365), .Z(n811) );
  ND2 U63 ( .A(n224), .B(n225), .Z(n1367) );
  ND2 U64 ( .A(n223), .B(n224), .Z(n1366) );
  ND2 U65 ( .A(n223), .B(n225), .Z(n1365) );
  ND3 U66 ( .A(n224), .B(n225), .C(n223), .Z(n788) );
  ND3 U67 ( .A(n279), .B(n277), .C(n278), .Z(n1880) );
  ND3 U68 ( .A(n613), .B(n277), .C(n278), .Z(n1958) );
  ND2 U69 ( .A(n223), .B(n224), .Z(n613) );
  ND3 U70 ( .A(n224), .B(n225), .C(n223), .Z(n508) );
  ND3 U71 ( .A(n224), .B(n225), .C(n223), .Z(n353) );
  ND3 U72 ( .A(n224), .B(n225), .C(n223), .Z(n335) );
  ND3 U73 ( .A(n2010), .B(n2009), .C(n2008), .Z(n307) );
  ND2 U74 ( .A(n278), .B(n277), .Z(n2010) );
  ND2 U75 ( .A(n306), .B(n278), .Z(n2009) );
  ND2 U76 ( .A(n278), .B(n279), .Z(n2008) );
  ND2 U77 ( .A(n224), .B(n225), .Z(n1440) );
  ND2 U78 ( .A(n223), .B(n224), .Z(n1009) );
  ND2 U79 ( .A(n223), .B(n224), .Z(n962) );
  ND2 U80 ( .A(n223), .B(n225), .Z(n1544) );
  ND2 U81 ( .A(n278), .B(n279), .Z(n2005) );
  ND2 U82 ( .A(n223), .B(n225), .Z(n1804) );
  ND2 U83 ( .A(n224), .B(n225), .Z(n1568) );
  ND2 U84 ( .A(n224), .B(n225), .Z(n1383) );
  ND2 U85 ( .A(n224), .B(n225), .Z(n1073) );
  ND2 U86 ( .A(n224), .B(n225), .Z(n996) );
  ND2 U87 ( .A(n223), .B(n224), .Z(n864) );
  ND2 U88 ( .A(n223), .B(n224), .Z(n733) );
  ND2 U89 ( .A(n223), .B(n225), .Z(n626) );
  ND2 U90 ( .A(n223), .B(n224), .Z(n636) );
  ND2 U91 ( .A(n223), .B(n224), .Z(n633) );
  ND2 U92 ( .A(n223), .B(n224), .Z(n955) );
  ND2 U93 ( .A(n223), .B(n225), .Z(n1101) );
  ND2 U94 ( .A(n223), .B(n224), .Z(n345) );
  ND2 U95 ( .A(n278), .B(n279), .Z(n2063) );
  ND2 U96 ( .A(n278), .B(n277), .Z(n2064) );
  ND2 U97 ( .A(n224), .B(n225), .Z(n549) );
  ND2 U98 ( .A(n279), .B(n277), .Z(n2034) );
  ND3 U99 ( .A(n224), .B(n225), .C(n223), .Z(n318) );
  ND3 U100 ( .A(n1931), .B(n1930), .C(n1929), .Z(n295) );
  ND2 U101 ( .A(n278), .B(n277), .Z(n1931) );
  ND2 U102 ( .A(n294), .B(n278), .Z(n1930) );
  ND2 U103 ( .A(n278), .B(n279), .Z(n1929) );
  AO7 U104 ( .A(n2213), .B(n2064), .C(n2063), .Z(n293) );
  IVP U105 ( .A(n292), .Z(n2213) );
  MUX41 U106 ( .D0(n860), .D1(n844), .D2(n853), .D3(n835), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N27) );
  MUX41 U107 ( .D0(n890), .D1(n878), .D2(n882), .D3(n869), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N28) );
  ND3 U108 ( .A(n2019), .B(n2018), .C(n2017), .Z(n882) );
  MUX41 U109 ( .D0(n826), .D1(n810), .D2(n818), .D3(n801), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N26) );
  MUX41 U110 ( .D0(n795), .D1(n780), .D2(n789), .D3(n772), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N25) );
  MUX41 U111 ( .D0(n737), .D1(n723), .D2(n729), .D3(n717), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N23) );
  MUX41 U112 ( .D0(n766), .D1(n749), .D2(n757), .D3(n745), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N24) );
  AO3 U113 ( .A(input_log2[43]), .B(n2096), .C(n278), .D(n2095), .Z(n566) );
  ND2 U114 ( .A(n1918), .B(n1917), .Z(N15) );
  ND2 U115 ( .A(input_log2[46]), .B(n220), .Z(n1918) );
  ND2 U116 ( .A(n570), .B(n220), .Z(n1917) );
  ND2 U117 ( .A(n2130), .B(n220), .Z(N16) );
  MUX21L U118 ( .A(n578), .B(n572), .S(input_log2[46]), .Z(n2130) );
  ND4 U119 ( .A(n2047), .B(n2046), .C(n2045), .D(n2044), .Z(n578) );
  ND2 U120 ( .A(n1916), .B(n1915), .Z(N17) );
  MUX21L U121 ( .A(n1914), .B(n1913), .S(input_log2[47]), .Z(n1916) );
  ND3 U122 ( .A(n581), .B(n220), .C(input_log2[46]), .Z(n1915) );
  MUX41 U123 ( .D0(n607), .D1(n594), .D2(n598), .D3(n592), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N18) );
  ND2 U124 ( .A(n1965), .B(n1964), .Z(n594) );
  ND2 U125 ( .A(n1881), .B(n1880), .Z(n592) );
  MUX41 U126 ( .D0(n629), .D1(n615), .D2(n621), .D3(n609), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N19) );
  ND2 U127 ( .A(n1879), .B(n1878), .Z(n609) );
  MUX41 U128 ( .D0(n653), .D1(n638), .D2(n645), .D3(n632), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N20) );
  ND3 U129 ( .A(n1875), .B(n1874), .C(n1873), .Z(n632) );
  MUX41 U130 ( .D0(n680), .D1(n666), .D2(n673), .D3(n658), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N21) );
  MUX41 U131 ( .D0(n709), .D1(n695), .D2(n701), .D3(n688), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N22) );
  MUX41 U132 ( .D0(n924), .D1(n907), .D2(n915), .D3(n898), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N29) );
  AO4 U133 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n631) );
  AO7 U134 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n571) );
  AO7 U135 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n292) );
  NR3 U136 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n582) );
  NR3 U137 ( .A(input_log2[43]), .B(n240), .C(input_log2[45]), .Z(n2050) );
  ND2 U138 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1751) );
  EO U139 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n276) );
  NR3 U140 ( .A(n241), .B(input_log2[43]), .C(input_log2[44]), .Z(n1852) );
  ND2 U141 ( .A(input_log2[42]), .B(n224), .Z(n1111) );
  NR3 U142 ( .A(n2210), .B(input_log2[44]), .C(input_log2[45]), .Z(n1848) );
  IVP U143 ( .A(n800), .Z(n2210) );
  AO7 U144 ( .A(input_log2[40]), .B(input_log2[41]), .C(n223), .Z(n800) );
  NR3 U145 ( .A(n242), .B(input_log2[44]), .C(input_log2[45]), .Z(n2106) );
  MUX21L U146 ( .A(n1117), .B(input_log2[42]), .S(input_log2[40]), .Z(n1120)
         );
  NR3 U147 ( .A(input_log2[45]), .B(input_log2[43]), .C(n2209), .Z(n1937) );
  IVP U148 ( .A(n779), .Z(n2209) );
  AO7 U149 ( .A(input_log2[41]), .B(n223), .C(n1360), .Z(n779) );
  ND2 U150 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1360) );
  NR3 U151 ( .A(n243), .B(input_log2[44]), .C(input_log2[45]), .Z(n2182) );
  ND2 U152 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1558) );
  NR3 U153 ( .A(input_log2[43]), .B(n1361), .C(input_log2[44]), .Z(n2136) );
  ND2 U154 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1361) );
  NR3 U155 ( .A(input_log2[42]), .B(input_log2[43]), .C(input_log2[45]), .Z(
        n1989) );
  NR3 U156 ( .A(n2207), .B(input_log2[43]), .C(input_log2[44]), .Z(n1984) );
  IVP U157 ( .A(n620), .Z(n2207) );
  AO7 U158 ( .A(input_log2[40]), .B(n223), .C(input_log2[41]), .Z(n620) );
  NR3 U159 ( .A(n244), .B(input_log2[44]), .C(input_log2[45]), .Z(n1980) );
  ND2 U160 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1539) );
  NR3 U161 ( .A(n245), .B(input_log2[43]), .C(input_log2[44]), .Z(n1862) );
  ND2 U162 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1143) );
  NR3 U163 ( .A(n246), .B(input_log2[44]), .C(input_log2[45]), .Z(n1858) );
  ND2 U164 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1104) );
  NR3 U165 ( .A(n247), .B(input_log2[43]), .C(input_log2[44]), .Z(n2197) );
  ND2 U166 ( .A(input_log2[42]), .B(n225), .Z(n1441) );
  NR3 U167 ( .A(input_log2[45]), .B(input_log2[44]), .C(n2206), .Z(n2194) );
  IVP U168 ( .A(n700), .Z(n2206) );
  AO7 U169 ( .A(input_log2[41]), .B(n223), .C(n1566), .Z(n700) );
  ND2 U170 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1566) );
  NR3 U171 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n803) );
  NR3 U172 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n647) );
  NR3 U173 ( .A(input_log2[45]), .B(input_log2[44]), .C(n248), .Z(n2087) );
  NR3 U174 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n301) );
  NR3 U175 ( .A(n249), .B(input_log2[43]), .C(input_log2[44]), .Z(n1887) );
  MUX21L U176 ( .A(n1122), .B(n1123), .S(input_log2[40]), .Z(n1127) );
  NR3 U177 ( .A(n225), .B(input_log2[44]), .C(input_log2[45]), .Z(n1883) );
  NR3 U178 ( .A(n250), .B(input_log2[44]), .C(input_log2[45]), .Z(n2118) );
  ND2 U179 ( .A(input_log2[42]), .B(input_log2[40]), .Z(n1130) );
  NR3 U180 ( .A(n251), .B(input_log2[43]), .C(input_log2[44]), .Z(n1974) );
  ND2 U181 ( .A(n224), .B(n225), .Z(n1228) );
  NR3 U182 ( .A(n252), .B(input_log2[43]), .C(input_log2[44]), .Z(n1897) );
  ND2 U183 ( .A(n223), .B(n224), .Z(n1140) );
  NR3 U184 ( .A(n253), .B(input_log2[44]), .C(input_log2[45]), .Z(n1893) );
  NR3 U185 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n478) );
  MUX41 U186 ( .D0(n958), .D1(n940), .D2(n949), .D3(n933), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N30) );
  AO4 U187 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n827) );
  AO7 U188 ( .A(input_log2[40]), .B(n224), .C(input_log2[42]), .Z(n834) );
  AO7 U189 ( .A(input_log2[42]), .B(n225), .C(n224), .Z(n840) );
  AO7 U190 ( .A(input_log2[40]), .B(input_log2[42]), .C(input_log2[41]), .Z(
        n851) );
  AO7 U191 ( .A(input_log2[41]), .B(n225), .C(input_log2[42]), .Z(n868) );
  AO7 U192 ( .A(input_log2[40]), .B(n223), .C(n224), .Z(n875) );
  AO7 U193 ( .A(input_log2[42]), .B(n224), .C(n225), .Z(n812) );
  AO7 U194 ( .A(input_log2[42]), .B(n224), .C(n1503), .Z(n815) );
  ND2 U195 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1503) );
  AO7 U196 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n819) );
  AO2 U197 ( .A(n2159), .B(n278), .C(n2158), .D(n720), .Z(n2167) );
  ND2 U198 ( .A(n1235), .B(n1234), .Z(n720) );
  NR2 U199 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2159) );
  NR2 U200 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2158) );
  AO4 U201 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[41]), .Z(n730) );
  AO2 U202 ( .A(n2135), .B(input_log2[44]), .C(n2134), .D(input_log2[44]), .Z(
        n2143) );
  NR2 U203 ( .A(input_log2[43]), .B(input_log2[40]), .Z(n2135) );
  NR2 U204 ( .A(input_log2[43]), .B(n278), .Z(n2134) );
  AO7 U205 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n758) );
  AO7 U206 ( .A(input_log2[40]), .B(n223), .C(n1792), .Z(n764) );
  ND2 U207 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1792) );
  AO3 U208 ( .A(n254), .B(n2005), .C(n2004), .D(n2003), .Z(n581) );
  MUX21L U209 ( .A(n2000), .B(n1999), .S(input_log2[44]), .Z(n2004) );
  MUX21L U210 ( .A(n2001), .B(n2002), .S(input_log2[43]), .Z(n2003) );
  AO7 U211 ( .A(input_log2[40]), .B(n224), .C(n223), .Z(n604) );
  AO7 U212 ( .A(input_log2[42]), .B(n224), .C(input_log2[40]), .Z(n652) );
  AO7 U213 ( .A(input_log2[42]), .B(n224), .C(n1164), .Z(n689) );
  ND2 U214 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1164) );
  AO2 U215 ( .A(n2147), .B(input_log2[45]), .C(n2146), .D(n939), .Z(n2155) );
  MUX21L U216 ( .A(input_log2[41]), .B(input_log2[40]), .S(input_log2[42]), 
        .Z(n939) );
  NR2 U217 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2147) );
  NR2 U218 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2146) );
  AO7 U219 ( .A(input_log2[40]), .B(n224), .C(input_log2[42]), .Z(n931) );
  AO7 U220 ( .A(input_log2[40]), .B(n223), .C(n1064), .Z(n894) );
  ND2 U221 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1064) );
  AO7 U222 ( .A(input_log2[40]), .B(n223), .C(n979), .Z(n891) );
  ND2 U223 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n979) );
  AO4 U224 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n904) );
  AO7 U225 ( .A(input_log2[41]), .B(n223), .C(n1203), .Z(n901) );
  ND2 U226 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1203) );
  AO7 U227 ( .A(input_log2[41]), .B(n223), .C(n1359), .Z(n906) );
  ND2 U228 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1359) );
  AO4 U229 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n294) );
  AO4 U230 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[41]), .Z(n547) );
  AO2 U231 ( .A(n2171), .B(n278), .C(n2170), .D(n505), .Z(n2179) );
  ND2 U232 ( .A(n1243), .B(n1242), .Z(n505) );
  NR2 U233 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2171) );
  NR2 U234 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2170) );
  AO7 U235 ( .A(input_log2[41]), .B(n223), .C(n1570), .Z(n515) );
  ND2 U236 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1570) );
  AO7 U237 ( .A(input_log2[40]), .B(n223), .C(input_log2[41]), .Z(n480) );
  AO7 U238 ( .A(input_log2[42]), .B(n225), .C(n1746), .Z(n492) );
  ND2 U239 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1746) );
  AO7 U240 ( .A(input_log2[42]), .B(n224), .C(input_log2[40]), .Z(n494) );
  AO4 U241 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n456) );
  AO7 U242 ( .A(input_log2[41]), .B(n223), .C(n1681), .Z(n459) );
  ND2 U243 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1681) );
  AO7 U244 ( .A(input_log2[40]), .B(input_log2[41]), .C(n223), .Z(n405) );
  AO7 U245 ( .A(input_log2[42]), .B(n224), .C(n1310), .Z(n414) );
  ND2 U246 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1310) );
  AO7 U247 ( .A(input_log2[40]), .B(n223), .C(n1793), .Z(n430) );
  ND2 U248 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1793) );
  AO7 U249 ( .A(input_log2[42]), .B(n225), .C(n224), .Z(n390) );
  AO4 U250 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n377) );
  AO7 U251 ( .A(input_log2[41]), .B(input_log2[42]), .C(n225), .Z(n396) );
  AO2 U252 ( .A(n315), .B(input_log2[45]), .C(input_log2[45]), .D(n279), .Z(
        n2032) );
  NR3 U253 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n315) );
  AO7 U254 ( .A(n277), .B(n1967), .C(n278), .Z(n305) );
  ND2 U255 ( .A(input_log2[44]), .B(n304), .Z(n1967) );
  ND2 U256 ( .A(n1294), .B(n223), .Z(n304) );
  ND2 U257 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1294) );
  AO7 U258 ( .A(n277), .B(n1968), .C(n278), .Z(n300) );
  ND2 U259 ( .A(input_log2[44]), .B(n299), .Z(n1968) );
  ND2 U260 ( .A(n1295), .B(n223), .Z(n299) );
  ND2 U261 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1295) );
  AO3 U262 ( .A(n278), .B(n1907), .C(n1906), .D(n1905), .Z(n347) );
  MUX21L U263 ( .A(n1902), .B(n1903), .S(input_log2[44]), .Z(n1906) );
  MUX21L U264 ( .A(n1904), .B(n279), .S(input_log2[43]), .Z(n1905) );
  ND2 U265 ( .A(n345), .B(n279), .Z(n1907) );
  AO7 U266 ( .A(n277), .B(n1966), .C(n278), .Z(n314) );
  ND2 U267 ( .A(input_log2[44]), .B(n313), .Z(n1966) );
  ND2 U268 ( .A(n1293), .B(n223), .Z(n313) );
  ND2 U269 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1293) );
  NR2 U270 ( .A(input_log2[40]), .B(n224), .Z(n1448) );
  NR2 U271 ( .A(input_log2[42]), .B(n224), .Z(n1117) );
  NR2 U272 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1576) );
  NR2 U273 ( .A(input_log2[41]), .B(n225), .Z(n1578) );
  NR2 U274 ( .A(input_log2[40]), .B(n223), .Z(n1766) );
  NR2 U275 ( .A(input_log2[40]), .B(n223), .Z(n1635) );
  NR2 U276 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n990) );
  NR2 U277 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1035) );
  NR2 U278 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n982) );
  NR2 U279 ( .A(n1119), .B(n1118), .Z(n1121) );
  NR2 U280 ( .A(input_log2[41]), .B(n223), .Z(n1119) );
  NR2 U281 ( .A(input_log2[41]), .B(n225), .Z(n1118) );
  NR2 U282 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1278) );
  NR2 U283 ( .A(input_log2[41]), .B(n223), .Z(n1279) );
  NR2 U284 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1434) );
  NR2 U285 ( .A(input_log2[40]), .B(n224), .Z(n1436) );
  NR2 U286 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1254) );
  NR2 U287 ( .A(input_log2[40]), .B(n224), .Z(n1256) );
  NR2 U288 ( .A(input_log2[41]), .B(n225), .Z(n1808) );
  NR2 U289 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1729) );
  NR2 U290 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1487) );
  NR2 U291 ( .A(input_log2[41]), .B(n225), .Z(n1517) );
  NR2 U292 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1177) );
  NR2 U293 ( .A(input_log2[42]), .B(n224), .Z(n1178) );
  NR2 U294 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1683) );
  NR2 U295 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1685) );
  NR2 U296 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1189) );
  NR2 U297 ( .A(input_log2[40]), .B(n223), .Z(n1191) );
  NR2 U298 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1337) );
  NR2 U299 ( .A(input_log2[41]), .B(n223), .Z(n1338) );
  NR2 U300 ( .A(input_log2[42]), .B(n224), .Z(n1216) );
  NR2 U301 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1215) );
  NR2 U302 ( .A(input_log2[40]), .B(n223), .Z(n1214) );
  NR2 U303 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1347) );
  NR2 U304 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1349) );
  NR2 U305 ( .A(input_log2[40]), .B(n223), .Z(n1353) );
  NR2 U306 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1719) );
  NR2 U307 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1721) );
  NR2 U308 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1039) );
  NR2 U309 ( .A(input_log2[41]), .B(n225), .Z(n1052) );
  NR2 U310 ( .A(input_log2[41]), .B(n223), .Z(n1053) );
  NR2 U311 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2053) );
  AN2P U312 ( .A(n279), .B(n567), .Z(n2049) );
  AO4 U313 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n567) );
  NR2 U314 ( .A(input_log2[43]), .B(n255), .Z(n2051) );
  ND2 U315 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1843) );
  NR2 U316 ( .A(input_log2[45]), .B(n279), .Z(n2002) );
  NR2 U317 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n2001) );
  NR2 U318 ( .A(input_log2[45]), .B(n256), .Z(n1999) );
  ND2 U319 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1512) );
  AN2P U320 ( .A(n277), .B(n580), .Z(n2000) );
  ND2 U321 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n580) );
  NR2 U322 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1532) );
  NR2 U323 ( .A(input_log2[41]), .B(n223), .Z(n1533) );
  NR2 U324 ( .A(input_log2[41]), .B(n225), .Z(n1528) );
  NR2 U325 ( .A(input_log2[41]), .B(n223), .Z(n1529) );
  NR2 U326 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1259) );
  NR2 U327 ( .A(input_log2[40]), .B(n224), .Z(n1261) );
  NR2 U328 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1236) );
  NR2 U329 ( .A(input_log2[41]), .B(n223), .Z(n1237) );
  NR2 U330 ( .A(input_log2[40]), .B(n223), .Z(n1692) );
  NR2 U331 ( .A(input_log2[44]), .B(n257), .Z(n2163) );
  ND2 U332 ( .A(input_log2[42]), .B(n224), .Z(n1323) );
  AN2P U333 ( .A(n277), .B(n722), .Z(n2161) );
  EO U334 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n722) );
  NR2 U335 ( .A(input_log2[43]), .B(n258), .Z(n2137) );
  ND2 U336 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1244) );
  NR2 U337 ( .A(input_log2[44]), .B(n277), .Z(n1994) );
  NR2 U338 ( .A(input_log2[44]), .B(n259), .Z(n1992) );
  EN U339 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1521) );
  NR2 U340 ( .A(input_log2[43]), .B(n279), .Z(n1957) );
  AN2P U341 ( .A(n278), .B(n614), .Z(n1954) );
  NR3 U342 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n614) );
  NR2 U343 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n1952) );
  NR2 U344 ( .A(input_log2[45]), .B(n279), .Z(n2195) );
  NR2 U345 ( .A(input_log2[41]), .B(n223), .Z(n832) );
  NR2 U346 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n830) );
  NR2 U347 ( .A(input_log2[41]), .B(n223), .Z(n839) );
  NR2 U348 ( .A(input_log2[41]), .B(n223), .Z(n887) );
  NR2 U349 ( .A(input_log2[42]), .B(n225), .Z(n888) );
  NR2 U350 ( .A(input_log2[40]), .B(n224), .Z(n814) );
  NR2 U351 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n750) );
  NR2 U352 ( .A(input_log2[40]), .B(n223), .Z(n754) );
  NR2 U353 ( .A(input_log2[40]), .B(n224), .Z(n756) );
  NR2 U354 ( .A(input_log2[46]), .B(n260), .Z(n1913) );
  ND2 U355 ( .A(n279), .B(n277), .Z(n1923) );
  NR2 U356 ( .A(input_log2[46]), .B(n2215), .Z(n1914) );
  IVP U357 ( .A(n590), .Z(n2215) );
  MUX21L U358 ( .A(n225), .B(n223), .S(input_log2[41]), .Z(n588) );
  NR2 U359 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n634) );
  NR2 U360 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n649) );
  NR2 U361 ( .A(input_log2[41]), .B(n223), .Z(n677) );
  NR2 U362 ( .A(input_log2[41]), .B(n225), .Z(n1311) );
  NR2 U363 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1551) );
  NR2 U364 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1004) );
  NR2 U365 ( .A(input_log2[41]), .B(n223), .Z(n1005) );
  NR2 U366 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1015) );
  NR2 U367 ( .A(input_log2[40]), .B(n224), .Z(n1017) );
  AN2P U368 ( .A(n279), .B(n935), .Z(n2150) );
  AO7 U369 ( .A(input_log2[41]), .B(n223), .C(n225), .Z(n935) );
  NR2 U370 ( .A(input_log2[43]), .B(n261), .Z(n2148) );
  ND2 U371 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1188) );
  NR2 U372 ( .A(input_log2[40]), .B(n223), .Z(n1315) );
  NR2 U373 ( .A(input_log2[42]), .B(n224), .Z(n908) );
  NR2 U374 ( .A(input_log2[40]), .B(n224), .Z(n910) );
  NR2 U375 ( .A(input_log2[41]), .B(n223), .Z(n1122) );
  NR2 U376 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1821) );
  NR2 U377 ( .A(input_log2[41]), .B(n225), .Z(n1823) );
  NR2 U378 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n998) );
  NR2 U379 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1056) );
  NR2 U380 ( .A(input_log2[41]), .B(n223), .Z(n1057) );
  NR2 U381 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1152) );
  NR2 U382 ( .A(input_log2[45]), .B(n279), .Z(n2088) );
  AN2P U383 ( .A(n278), .B(n311), .Z(n2086) );
  AO7 U384 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n311) );
  NR2 U385 ( .A(input_log2[40]), .B(n223), .Z(n1560) );
  NR2 U386 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1702) );
  NR2 U387 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1834) );
  NR2 U388 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1835) );
  NR2 U389 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1620) );
  NR2 U390 ( .A(input_log2[41]), .B(n223), .Z(n1621) );
  NR2 U391 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1086) );
  NR2 U392 ( .A(input_log2[40]), .B(n224), .Z(n1088) );
  NR2 U393 ( .A(input_log2[42]), .B(n224), .Z(n1198) );
  NR2 U394 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1197) );
  NR2 U395 ( .A(input_log2[40]), .B(n223), .Z(n1196) );
  NR2 U396 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1172) );
  NR2 U397 ( .A(input_log2[40]), .B(n224), .Z(n1174) );
  NR2 U398 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1230) );
  NR2 U399 ( .A(input_log2[41]), .B(n225), .Z(n1455) );
  NR2 U400 ( .A(input_log2[41]), .B(n223), .Z(n1456) );
  NR2 U401 ( .A(input_log2[40]), .B(n224), .Z(n1627) );
  NR2 U402 ( .A(input_log2[40]), .B(n223), .Z(n1628) );
  NR2 U403 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1736) );
  NR2 U404 ( .A(input_log2[41]), .B(n225), .Z(n1738) );
  AN2P U405 ( .A(n277), .B(n297), .Z(n2103) );
  AO4 U406 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n297) );
  NR2 U407 ( .A(n1133), .B(n1132), .Z(n1135) );
  NR2 U408 ( .A(input_log2[41]), .B(n223), .Z(n1133) );
  NR2 U409 ( .A(input_log2[41]), .B(n225), .Z(n1132) );
  AN2P U410 ( .A(n278), .B(n346), .Z(n1902) );
  AN3 U411 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .Z(
        n346) );
  NR2 U412 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2025) );
  AN2P U413 ( .A(n279), .B(n330), .Z(n2021) );
  AO4 U414 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n330) );
  NR2 U415 ( .A(input_log2[41]), .B(n225), .Z(n548) );
  NR2 U416 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n524) );
  NR2 U417 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n463) );
  NR2 U418 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n354) );
  NR2 U419 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n336) );
  NR2 U420 ( .A(n1910), .B(n1909), .Z(n1912) );
  NR2 U421 ( .A(input_log2[45]), .B(n277), .Z(n1910) );
  NR2 U422 ( .A(input_log2[45]), .B(n262), .Z(n1909) );
  NR2 U423 ( .A(n1926), .B(n1925), .Z(n1928) );
  NR2 U424 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n1926) );
  NR2 U425 ( .A(input_log2[44]), .B(n263), .Z(n1925) );
  ND2 U426 ( .A(n1815), .B(n1814), .Z(n557) );
  ND2 U427 ( .A(n223), .B(n225), .Z(n1815) );
  ND2 U428 ( .A(input_log2[41]), .B(n223), .Z(n1814) );
  ND3 U429 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n558) );
  NR2 U430 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n556) );
  ND3 U431 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .Z(
        n312) );
  MUX21L U432 ( .A(n224), .B(n1811), .S(input_log2[40]), .Z(n1813) );
  ND2 U433 ( .A(input_log2[42]), .B(n224), .Z(n1812) );
  NR2 U434 ( .A(input_log2[42]), .B(n224), .Z(n1811) );
  ND2 U435 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1574) );
  EO U436 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1575) );
  ND4 U437 ( .A(n577), .B(input_log2[44]), .C(n278), .D(n277), .Z(n2044) );
  ND2 U438 ( .A(n1731), .B(n1730), .Z(n577) );
  MUX21L U439 ( .A(n1728), .B(n225), .S(input_log2[41]), .Z(n1730) );
  AO6 U440 ( .A(input_log2[41]), .B(n223), .C(n1729), .Z(n1731) );
  ND4 U441 ( .A(n858), .B(input_log2[44]), .C(n278), .D(n277), .Z(n2071) );
  AO7 U442 ( .A(input_log2[41]), .B(n225), .C(n223), .Z(n858) );
  ND4 U443 ( .A(n799), .B(input_log2[44]), .C(n278), .D(n277), .Z(n1853) );
  ND2 U444 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n799) );
  ND4 U445 ( .A(n777), .B(input_log2[44]), .C(n278), .D(n277), .Z(n1938) );
  MUX21L U446 ( .A(n1306), .B(n1305), .S(input_log2[40]), .Z(n777) );
  ND2 U447 ( .A(n223), .B(n224), .Z(n1306) );
  ND2 U448 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1305) );
  ND4 U449 ( .A(n619), .B(input_log2[44]), .C(n278), .D(n277), .Z(n1985) );
  ND2 U450 ( .A(n1508), .B(n1507), .Z(n619) );
  ND2 U451 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1507) );
  EO U452 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1508) );
  ND4 U453 ( .A(n657), .B(input_log2[44]), .C(n278), .D(n277), .Z(n1863) );
  NR2 U454 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n657) );
  ND4 U455 ( .A(n2074), .B(n2073), .C(n2072), .D(n2071), .Z(n860) );
  MUX21L U456 ( .A(n2065), .B(n2066), .S(input_log2[43]), .Z(n2074) );
  MUX21L U457 ( .A(n2067), .B(n2068), .S(input_log2[44]), .Z(n2073) );
  MUX21L U458 ( .A(n2070), .B(n2069), .S(input_log2[44]), .Z(n2072) );
  ND4 U459 ( .A(n1856), .B(n1855), .C(n1854), .D(n1853), .Z(n801) );
  MUX21L U460 ( .A(n1847), .B(n1848), .S(input_log2[43]), .Z(n1856) );
  MUX21L U461 ( .A(n1849), .B(n1850), .S(input_log2[43]), .Z(n1855) );
  MUX21L U462 ( .A(n1852), .B(n1851), .S(input_log2[45]), .Z(n1854) );
  ND4 U463 ( .A(n2117), .B(n2116), .C(n2115), .D(n2114), .Z(n772) );
  MUX21L U464 ( .A(n2106), .B(n2107), .S(input_log2[43]), .Z(n2117) );
  MUX21L U465 ( .A(n2108), .B(n2109), .S(input_log2[45]), .Z(n2116) );
  MUX21L U466 ( .A(n2110), .B(n2111), .S(input_log2[43]), .Z(n2115) );
  ND4 U467 ( .A(n1941), .B(n1940), .C(n1939), .D(n1938), .Z(n780) );
  MUX21L U468 ( .A(n1932), .B(n1933), .S(input_log2[43]), .Z(n1941) );
  MUX21L U469 ( .A(n1934), .B(n1935), .S(input_log2[44]), .Z(n1940) );
  MUX21L U470 ( .A(n1937), .B(n1936), .S(input_log2[44]), .Z(n1939) );
  ND4 U471 ( .A(n2169), .B(n2168), .C(n2167), .D(n2166), .Z(n723) );
  MUX21L U472 ( .A(n2161), .B(n2160), .S(input_log2[45]), .Z(n2169) );
  MUX21L U473 ( .A(n2163), .B(n2162), .S(input_log2[45]), .Z(n2168) );
  MUX21L U474 ( .A(n2165), .B(n2164), .S(input_log2[45]), .Z(n2166) );
  ND4 U475 ( .A(n2193), .B(n2192), .C(n2191), .D(n2190), .Z(n729) );
  MUX21L U476 ( .A(n2182), .B(n2183), .S(input_log2[43]), .Z(n2193) );
  MUX21L U477 ( .A(n2184), .B(n2185), .S(input_log2[45]), .Z(n2192) );
  MUX21L U478 ( .A(n2186), .B(n2187), .S(input_log2[43]), .Z(n2191) );
  ND4 U479 ( .A(n2145), .B(n2144), .C(n2143), .D(n2142), .Z(n749) );
  MUX21L U480 ( .A(n2136), .B(n2137), .S(input_log2[45]), .Z(n2145) );
  MUX21L U481 ( .A(n2139), .B(n2138), .S(input_log2[45]), .Z(n2144) );
  MUX21L U482 ( .A(n2141), .B(n2140), .S(input_log2[45]), .Z(n2142) );
  ND4 U483 ( .A(n1998), .B(n1997), .C(n1996), .D(n1995), .Z(n598) );
  MUX21L U484 ( .A(n1989), .B(n1990), .S(input_log2[44]), .Z(n1998) );
  MUX21L U485 ( .A(n1991), .B(n1992), .S(input_log2[43]), .Z(n1997) );
  MUX21L U486 ( .A(n1993), .B(n1994), .S(input_log2[45]), .Z(n1996) );
  ND4 U487 ( .A(n1961), .B(n1960), .C(n1959), .D(n1958), .Z(n615) );
  MUX21L U488 ( .A(n1952), .B(n1953), .S(input_log2[43]), .Z(n1961) );
  MUX21L U489 ( .A(n1954), .B(n1955), .S(input_log2[44]), .Z(n1960) );
  MUX21L U490 ( .A(n1956), .B(n1957), .S(input_log2[45]), .Z(n1959) );
  ND4 U491 ( .A(n1988), .B(n1987), .C(n1986), .D(n1985), .Z(n621) );
  MUX21L U492 ( .A(n1979), .B(n1980), .S(input_log2[43]), .Z(n1988) );
  MUX21L U493 ( .A(n1981), .B(n1982), .S(input_log2[43]), .Z(n1987) );
  MUX21L U494 ( .A(n1984), .B(n1983), .S(input_log2[45]), .Z(n1986) );
  ND4 U495 ( .A(n1866), .B(n1865), .C(n1864), .D(n1863), .Z(n658) );
  MUX21L U496 ( .A(n1857), .B(n1858), .S(input_log2[43]), .Z(n1866) );
  MUX21L U497 ( .A(n1859), .B(n1860), .S(input_log2[43]), .Z(n1865) );
  MUX21L U498 ( .A(n1862), .B(n1861), .S(input_log2[45]), .Z(n1864) );
  ND4 U499 ( .A(n2205), .B(n2204), .C(n2203), .D(n2202), .Z(n701) );
  MUX21L U500 ( .A(n2194), .B(n2195), .S(input_log2[43]), .Z(n2205) );
  MUX21L U501 ( .A(n2196), .B(n2197), .S(input_log2[45]), .Z(n2204) );
  MUX21L U502 ( .A(n2198), .B(n2199), .S(input_log2[45]), .Z(n2203) );
  ND4 U503 ( .A(n2157), .B(n2156), .C(n2155), .D(n2154), .Z(n940) );
  MUX21L U504 ( .A(n2149), .B(n2148), .S(input_log2[45]), .Z(n2157) );
  MUX21L U505 ( .A(n2151), .B(n2150), .S(input_log2[45]), .Z(n2156) );
  MUX21L U506 ( .A(n2153), .B(n2152), .S(input_log2[45]), .Z(n2154) );
  ND4 U507 ( .A(n529), .B(input_log2[44]), .C(n278), .D(n277), .Z(n1888) );
  MUX21L U508 ( .A(n1074), .B(input_log2[40]), .S(input_log2[42]), .Z(n529) );
  ND2 U509 ( .A(input_log2[40]), .B(n224), .Z(n1074) );
  ND4 U510 ( .A(n473), .B(input_log2[44]), .C(input_log2[45]), .D(n277), .Z(
        n1975) );
  ND2 U511 ( .A(n1183), .B(n1182), .Z(n473) );
  ND2 U512 ( .A(n223), .B(n224), .Z(n1182) );
  EO U513 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1183) );
  ND4 U514 ( .A(input_log2[42]), .B(input_log2[44]), .C(n278), .D(n277), .Z(
        n1898) );
  ND4 U515 ( .A(n322), .B(input_log2[44]), .C(n278), .D(n277), .Z(n2081) );
  ND2 U516 ( .A(n1756), .B(n1755), .Z(n322) );
  ND2 U517 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1756) );
  ND2 U518 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1755) );
  ND4 U519 ( .A(n1891), .B(n1890), .C(n1889), .D(n1888), .Z(n530) );
  MUX21L U520 ( .A(n1882), .B(n1883), .S(input_log2[43]), .Z(n1891) );
  MUX21L U521 ( .A(n1884), .B(n1885), .S(input_log2[43]), .Z(n1890) );
  MUX21L U522 ( .A(n1887), .B(n1886), .S(input_log2[45]), .Z(n1889) );
  ND4 U523 ( .A(n2129), .B(n2128), .C(n2127), .D(n2126), .Z(n502) );
  MUX21L U524 ( .A(n2118), .B(n2119), .S(input_log2[43]), .Z(n2129) );
  MUX21L U525 ( .A(n2120), .B(n2121), .S(input_log2[45]), .Z(n2128) );
  MUX21L U526 ( .A(n2122), .B(n2123), .S(input_log2[43]), .Z(n2127) );
  ND4 U527 ( .A(n1978), .B(n1977), .C(n1976), .D(n1975), .Z(n477) );
  MUX21L U528 ( .A(n1969), .B(n1970), .S(input_log2[43]), .Z(n1978) );
  MUX21L U529 ( .A(n1971), .B(n1972), .S(input_log2[44]), .Z(n1977) );
  MUX21L U530 ( .A(n1973), .B(n1974), .S(input_log2[45]), .Z(n1976) );
  ND4 U531 ( .A(n1901), .B(n1900), .C(n1899), .D(n1898), .Z(n374) );
  MUX21L U532 ( .A(n1892), .B(n1893), .S(input_log2[43]), .Z(n1901) );
  MUX21L U533 ( .A(n1894), .B(n1895), .S(input_log2[43]), .Z(n1900) );
  MUX21L U534 ( .A(n1897), .B(n1896), .S(input_log2[45]), .Z(n1899) );
  ND4 U535 ( .A(n2029), .B(n2028), .C(n2027), .D(n2026), .Z(n334) );
  MUX21L U536 ( .A(n2020), .B(n2021), .S(input_log2[45]), .Z(n2029) );
  MUX21L U537 ( .A(n2022), .B(n2023), .S(input_log2[44]), .Z(n2028) );
  MUX21L U538 ( .A(n2024), .B(n2025), .S(input_log2[45]), .Z(n2027) );
  ND2 U539 ( .A(n1082), .B(n1081), .Z(n833) );
  ND2 U540 ( .A(n1010), .B(n1009), .Z(n829) );
  ND2 U541 ( .A(n1050), .B(n1049), .Z(n831) );
  MUX21L U542 ( .A(n988), .B(input_log2[41]), .S(input_log2[42]), .Z(n863) );
  MUX21L U543 ( .A(n964), .B(n963), .S(input_log2[41]), .Z(n862) );
  MUX21L U544 ( .A(n962), .B(n961), .S(input_log2[40]), .Z(n861) );
  MUX21L U545 ( .A(n1614), .B(n225), .S(input_log2[41]), .Z(n884) );
  ND2 U546 ( .A(n1800), .B(n1799), .Z(n889) );
  MUX21L U547 ( .A(n1556), .B(input_log2[41]), .S(input_log2[42]), .Z(n817) );
  MUX21L U548 ( .A(n1414), .B(n1413), .S(input_log2[40]), .Z(n813) );
  MUX21L U549 ( .A(n1544), .B(n223), .S(input_log2[41]), .Z(n816) );
  MUX21L U550 ( .A(input_log2[42]), .B(input_log2[41]), .S(input_log2[40]), 
        .Z(n755) );
  ND2 U551 ( .A(n1466), .B(n1465), .Z(n753) );
  MUX21L U552 ( .A(n1804), .B(n1803), .S(input_log2[41]), .Z(n606) );
  ND2 U553 ( .A(n1699), .B(n1698), .Z(n603) );
  ND2 U554 ( .A(n1609), .B(n1608), .Z(n600) );
  ND2 U555 ( .A(n1328), .B(n1327), .Z(n637) );
  ND2 U556 ( .A(n1210), .B(n223), .Z(n635) );
  MUX21L U557 ( .A(n224), .B(n1383), .S(input_log2[42]), .Z(n639) );
  ND2 U558 ( .A(n1569), .B(n1568), .Z(n644) );
  ND2 U559 ( .A(n1492), .B(n1491), .Z(n642) );
  MUX21L U560 ( .A(n224), .B(n1382), .S(input_log2[40]), .Z(n667) );
  ND2 U561 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n672) );
  ND2 U562 ( .A(n1421), .B(n1420), .Z(n668) );
  MUX21L U563 ( .A(input_log2[41]), .B(n1116), .S(input_log2[40]), .Z(n687) );
  MUX21L U564 ( .A(n224), .B(n996), .S(input_log2[42]), .Z(n682) );
  MUX21L U565 ( .A(n224), .B(n1073), .S(input_log2[42]), .Z(n685) );
  MUX21L U566 ( .A(n1110), .B(n1109), .S(input_log2[42]), .Z(n897) );
  MUX21L U567 ( .A(input_log2[42]), .B(n1024), .S(input_log2[40]), .Z(n893) );
  MUX21L U568 ( .A(n223), .B(n224), .S(input_log2[40]), .Z(n895) );
  MUX21L U569 ( .A(n225), .B(n224), .S(input_log2[42]), .Z(n913) );
  MUX21L U570 ( .A(input_log2[42]), .B(n1469), .S(input_log2[40]), .Z(n912) );
  ND2 U571 ( .A(n1135), .B(n1134), .Z(n439) );
  ND2 U572 ( .A(n1023), .B(n1022), .Z(n435) );
  ND2 U573 ( .A(n1079), .B(n1078), .Z(n437) );
  ND2 U574 ( .A(n1102), .B(n1101), .Z(n406) );
  ND2 U575 ( .A(n1003), .B(n1002), .Z(n402) );
  ND2 U576 ( .A(n1047), .B(n1046), .Z(n404) );
  EO U577 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1752) );
  EO U578 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1844) );
  EN U579 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1245) );
  EN U580 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1520) );
  AN3 U581 ( .A(input_log2[44]), .B(n568), .C(input_log2[43]), .Z(n2052) );
  NR2 U582 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n568) );
  AN3 U583 ( .A(n569), .B(n279), .C(input_log2[43]), .Z(n2048) );
  ND3 U584 ( .A(n1778), .B(n1777), .C(n1776), .Z(n569) );
  ND2 U585 ( .A(input_log2[40]), .B(n224), .Z(n1778) );
  ND2 U586 ( .A(n223), .B(n224), .Z(n1777) );
  AN3 U587 ( .A(n857), .B(n278), .C(input_log2[43]), .Z(n2069) );
  MUX21L U588 ( .A(n223), .B(n224), .S(input_log2[40]), .Z(n857) );
  AN3 U589 ( .A(n854), .B(input_log2[43]), .C(input_log2[45]), .Z(n2068) );
  ND2 U590 ( .A(n1580), .B(n1579), .Z(n854) );
  MUX21L U591 ( .A(n1577), .B(n1578), .S(input_log2[42]), .Z(n1580) );
  ND2 U592 ( .A(n1576), .B(n224), .Z(n1579) );
  AN3 U593 ( .A(n859), .B(n278), .C(input_log2[43]), .Z(n2067) );
  ND2 U594 ( .A(n1768), .B(n1767), .Z(n859) );
  MUX21L U595 ( .A(n1765), .B(n1766), .S(input_log2[41]), .Z(n1768) );
  ND3 U596 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1767) );
  AN3 U597 ( .A(n855), .B(n279), .C(input_log2[45]), .Z(n2066) );
  ND2 U598 ( .A(n1637), .B(n1636), .Z(n855) );
  MUX21L U599 ( .A(n1634), .B(n1635), .S(input_log2[41]), .Z(n1637) );
  ND3 U600 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1636) );
  AN3 U601 ( .A(n856), .B(n279), .C(input_log2[45]), .Z(n2065) );
  ND2 U602 ( .A(input_log2[42]), .B(n225), .Z(n856) );
  EO U603 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1050) );
  EO U604 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1010) );
  AN3 U605 ( .A(n797), .B(n279), .C(input_log2[43]), .Z(n1851) );
  ND2 U606 ( .A(n992), .B(n991), .Z(n797) );
  MUX21L U607 ( .A(n989), .B(n225), .S(input_log2[41]), .Z(n991) );
  AO6 U608 ( .A(input_log2[41]), .B(n223), .C(n990), .Z(n992) );
  AN3 U609 ( .A(n798), .B(n278), .C(input_log2[44]), .Z(n1850) );
  MUX21L U610 ( .A(n225), .B(n1033), .S(input_log2[41]), .Z(n798) );
  ND2 U611 ( .A(n223), .B(n225), .Z(n1033) );
  AN3 U612 ( .A(n796), .B(input_log2[45]), .C(input_log2[44]), .Z(n1849) );
  ND2 U613 ( .A(n981), .B(n980), .Z(n796) );
  ND2 U614 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n980) );
  EN U615 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n981) );
  AN3 U616 ( .A(n225), .B(n279), .C(input_log2[45]), .Z(n1847) );
  ND2 U617 ( .A(n1037), .B(n1036), .Z(n769) );
  MUX21L U618 ( .A(n1034), .B(n225), .S(input_log2[41]), .Z(n1036) );
  AO6 U619 ( .A(input_log2[41]), .B(n223), .C(n1035), .Z(n1037) );
  AN3 U620 ( .A(n224), .B(n279), .C(input_log2[45]), .Z(n2110) );
  ND2 U621 ( .A(n984), .B(n983), .Z(n767) );
  MUX21L U622 ( .A(n982), .B(input_log2[42]), .S(input_log2[40]), .Z(n984) );
  ND2 U623 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n983) );
  AN3 U624 ( .A(n770), .B(n277), .C(input_log2[44]), .Z(n2108) );
  ND2 U625 ( .A(n1069), .B(n1068), .Z(n770) );
  MUX21L U626 ( .A(n1067), .B(n223), .S(input_log2[40]), .Z(n1069) );
  ND2 U627 ( .A(input_log2[40]), .B(n224), .Z(n1068) );
  AN3 U628 ( .A(n776), .B(n278), .C(input_log2[43]), .Z(n1936) );
  ND2 U629 ( .A(n1277), .B(n1276), .Z(n776) );
  MUX21L U630 ( .A(n224), .B(n1275), .S(input_log2[42]), .Z(n1277) );
  ND2 U631 ( .A(n224), .B(n225), .Z(n1276) );
  AN3 U632 ( .A(n773), .B(input_log2[43]), .C(input_log2[45]), .Z(n1935) );
  MUX21L U633 ( .A(n1145), .B(input_log2[41]), .S(input_log2[42]), .Z(n773) );
  ND2 U634 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1145) );
  AN3 U635 ( .A(n778), .B(n278), .C(input_log2[43]), .Z(n1934) );
  MUX21L U636 ( .A(n225), .B(n224), .S(input_log2[42]), .Z(n778) );
  AN3 U637 ( .A(n774), .B(n279), .C(input_log2[45]), .Z(n1933) );
  AO7 U638 ( .A(input_log2[40]), .B(n223), .C(input_log2[41]), .Z(n774) );
  AN3 U639 ( .A(n775), .B(n279), .C(input_log2[45]), .Z(n1932) );
  ND2 U640 ( .A(n1221), .B(n1220), .Z(n775) );
  MUX21L U641 ( .A(n1219), .B(n223), .S(input_log2[40]), .Z(n1221) );
  ND2 U642 ( .A(input_log2[40]), .B(n224), .Z(n1220) );
  AN3 U643 ( .A(input_log2[43]), .B(input_log2[44]), .C(n718), .Z(n2164) );
  ND2 U644 ( .A(n1163), .B(n1162), .Z(n718) );
  MUX21L U645 ( .A(n225), .B(n1161), .S(input_log2[42]), .Z(n1163) );
  ND2 U646 ( .A(n224), .B(n225), .Z(n1162) );
  AN3 U647 ( .A(input_log2[44]), .B(n721), .C(input_log2[43]), .Z(n2165) );
  ND2 U648 ( .A(n1282), .B(n1281), .Z(n721) );
  MUX21L U649 ( .A(n1279), .B(n1280), .S(input_log2[40]), .Z(n1282) );
  ND2 U650 ( .A(n1278), .B(input_log2[40]), .Z(n1281) );
  AN3 U651 ( .A(n719), .B(n279), .C(input_log2[43]), .Z(n2162) );
  EO U652 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n719) );
  AN3 U653 ( .A(n225), .B(n277), .C(input_log2[44]), .Z(n2160) );
  NR2 U654 ( .A(n279), .B(n280), .Z(n2187) );
  ND3 U655 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .Z(
        n280) );
  AN3 U656 ( .A(n726), .B(n279), .C(input_log2[45]), .Z(n2186) );
  ND2 U657 ( .A(n1438), .B(n1437), .Z(n726) );
  MUX21L U658 ( .A(n1435), .B(n1436), .S(input_log2[42]), .Z(n1438) );
  ND2 U659 ( .A(n1434), .B(n225), .Z(n1437) );
  MUX21L U660 ( .A(input_log2[41]), .B(n1381), .S(input_log2[40]), .Z(n724) );
  ND2 U661 ( .A(input_log2[41]), .B(n223), .Z(n1381) );
  AN3 U662 ( .A(n727), .B(n277), .C(input_log2[44]), .Z(n2184) );
  MUX21L U663 ( .A(input_log2[40]), .B(input_log2[41]), .S(input_log2[42]), 
        .Z(n727) );
  ND2 U664 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n746) );
  AN3 U665 ( .A(input_log2[43]), .B(n747), .C(input_log2[44]), .Z(n2141) );
  ND2 U666 ( .A(n1258), .B(n1257), .Z(n747) );
  MUX21L U667 ( .A(n1255), .B(n1256), .S(input_log2[42]), .Z(n1258) );
  ND2 U668 ( .A(n1254), .B(n225), .Z(n1257) );
  AN3 U669 ( .A(input_log2[42]), .B(n279), .C(input_log2[43]), .Z(n2138) );
  AN3 U670 ( .A(n748), .B(n279), .C(input_log2[43]), .Z(n2139) );
  ND2 U671 ( .A(n1321), .B(n1320), .Z(n748) );
  MUX21L U672 ( .A(n1319), .B(n223), .S(input_log2[41]), .Z(n1321) );
  ND2 U673 ( .A(input_log2[41]), .B(n225), .Z(n1320) );
  EO U674 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1466) );
  AN3 U675 ( .A(n596), .B(input_log2[43]), .C(input_log2[44]), .Z(n1993) );
  AO7 U676 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n596) );
  AN3 U677 ( .A(n597), .B(n278), .C(input_log2[44]), .Z(n1991) );
  ND2 U678 ( .A(n1510), .B(n1509), .Z(n597) );
  ND2 U679 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1510) );
  ND2 U680 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1509) );
  AN3 U681 ( .A(n595), .B(n277), .C(input_log2[45]), .Z(n1990) );
  NR2 U682 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n595) );
  AN3 U683 ( .A(n612), .B(input_log2[43]), .C(input_log2[44]), .Z(n1956) );
  ND2 U684 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n612) );
  NR2 U685 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n610) );
  AN3 U686 ( .A(n611), .B(n279), .C(input_log2[45]), .Z(n1953) );
  ND2 U687 ( .A(n1211), .B(n223), .Z(n611) );
  ND2 U688 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1211) );
  AN3 U689 ( .A(n223), .B(n279), .C(input_log2[43]), .Z(n1983) );
  AN3 U690 ( .A(n618), .B(n278), .C(input_log2[44]), .Z(n1982) );
  ND2 U691 ( .A(n1489), .B(n1488), .Z(n618) );
  MUX21L U692 ( .A(n1487), .B(input_log2[42]), .S(input_log2[40]), .Z(n1489)
         );
  ND2 U693 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1488) );
  AN3 U694 ( .A(n616), .B(input_log2[45]), .C(input_log2[44]), .Z(n1981) );
  ND2 U695 ( .A(n223), .B(n224), .Z(n616) );
  AN3 U696 ( .A(n617), .B(n279), .C(input_log2[45]), .Z(n1979) );
  EN U697 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n617) );
  AN3 U698 ( .A(n655), .B(n279), .C(input_log2[43]), .Z(n1861) );
  NR2 U699 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n655) );
  AN3 U700 ( .A(n656), .B(n278), .C(input_log2[44]), .Z(n1860) );
  AO7 U701 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n656) );
  AN3 U702 ( .A(n654), .B(input_log2[45]), .C(input_log2[44]), .Z(n1859) );
  ND3 U703 ( .A(n224), .B(n225), .C(n223), .Z(n654) );
  AN3 U704 ( .A(input_log2[42]), .B(n279), .C(input_log2[45]), .Z(n1857) );
  AN3 U705 ( .A(n696), .B(n277), .C(input_log2[44]), .Z(n2199) );
  ND2 U706 ( .A(n1394), .B(n1393), .Z(n696) );
  ND2 U707 ( .A(input_log2[41]), .B(n223), .Z(n1393) );
  EO U708 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1394) );
  ND2 U709 ( .A(n1519), .B(n1518), .Z(n699) );
  MUX21L U710 ( .A(n225), .B(n1517), .S(input_log2[42]), .Z(n1519) );
  ND2 U711 ( .A(input_log2[41]), .B(n223), .Z(n1518) );
  ND2 U712 ( .A(input_log2[41]), .B(n223), .Z(n698) );
  EN U713 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n740) );
  EN U714 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n601) );
  EN U715 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n602) );
  EO U716 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n1964) );
  EO U717 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n623) );
  EO U718 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n641) );
  EN U719 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n670) );
  EO U720 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n660) );
  AN3 U721 ( .A(input_log2[43]), .B(input_log2[44]), .C(n934), .Z(n2152) );
  MUX21L U722 ( .A(input_log2[41]), .B(input_log2[40]), .S(input_log2[42]), 
        .Z(n934) );
  AN3 U723 ( .A(input_log2[44]), .B(n936), .C(input_log2[43]), .Z(n2153) );
  ND2 U724 ( .A(n223), .B(n225), .Z(n936) );
  AN3 U725 ( .A(n938), .B(n279), .C(input_log2[43]), .Z(n2151) );
  MUX21L U726 ( .A(n1336), .B(n225), .S(input_log2[41]), .Z(n938) );
  ND2 U727 ( .A(input_log2[42]), .B(n225), .Z(n1336) );
  AN3 U728 ( .A(n937), .B(n277), .C(input_log2[44]), .Z(n2149) );
  ND2 U729 ( .A(n1313), .B(n1312), .Z(n937) );
  MUX21L U730 ( .A(n1311), .B(n225), .S(input_log2[42]), .Z(n1313) );
  ND2 U731 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1312) );
  EO U732 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n902) );
  AN3 U733 ( .A(n309), .B(n279), .C(input_log2[45]), .Z(n2085) );
  AO4 U734 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n309) );
  ND2 U735 ( .A(n1760), .B(n1759), .Z(n302) );
  ND2 U736 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1760) );
  ND2 U737 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1759) );
  EO U738 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1797) );
  AN3 U739 ( .A(n527), .B(n279), .C(input_log2[43]), .Z(n1886) );
  ND2 U740 ( .A(n1000), .B(n999), .Z(n527) );
  MUX21L U741 ( .A(n997), .B(n225), .S(input_log2[42]), .Z(n999) );
  AO6 U742 ( .A(input_log2[42]), .B(n224), .C(n998), .Z(n1000) );
  AN3 U743 ( .A(n528), .B(n278), .C(input_log2[44]), .Z(n1885) );
  ND2 U744 ( .A(n1060), .B(n1059), .Z(n528) );
  MUX21L U745 ( .A(n1057), .B(n1058), .S(input_log2[40]), .Z(n1060) );
  ND2 U746 ( .A(n1056), .B(input_log2[40]), .Z(n1059) );
  AN3 U747 ( .A(n526), .B(input_log2[45]), .C(input_log2[44]), .Z(n1884) );
  ND2 U748 ( .A(n223), .B(n224), .Z(n526) );
  AN3 U749 ( .A(input_log2[41]), .B(n279), .C(input_log2[45]), .Z(n1882) );
  ND3 U750 ( .A(n1063), .B(n1062), .C(n1061), .Z(n499) );
  ND2 U751 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1063) );
  ND2 U752 ( .A(input_log2[40]), .B(n223), .Z(n1062) );
  AN3 U753 ( .A(n498), .B(n279), .C(input_log2[45]), .Z(n2122) );
  EN U754 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n498) );
  ND2 U755 ( .A(n223), .B(n224), .Z(n496) );
  AN3 U756 ( .A(n500), .B(n277), .C(input_log2[44]), .Z(n2120) );
  ND2 U757 ( .A(n1076), .B(n1075), .Z(n500) );
  ND2 U758 ( .A(n224), .B(n225), .Z(n1076) );
  ND2 U759 ( .A(input_log2[42]), .B(n224), .Z(n1075) );
  AN3 U760 ( .A(input_log2[44]), .B(n474), .C(input_log2[43]), .Z(n1973) );
  ND3 U761 ( .A(n1285), .B(n1284), .C(n1283), .Z(n474) );
  ND2 U762 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1285) );
  ND2 U763 ( .A(input_log2[40]), .B(n223), .Z(n1284) );
  AN3 U764 ( .A(input_log2[43]), .B(input_log2[45]), .C(n472), .Z(n1972) );
  ND2 U765 ( .A(n1154), .B(n1153), .Z(n472) );
  MUX21L U766 ( .A(n1151), .B(n225), .S(input_log2[41]), .Z(n1153) );
  AO6 U767 ( .A(input_log2[41]), .B(n223), .C(n1152), .Z(n1154) );
  AN3 U768 ( .A(n476), .B(n278), .C(input_log2[43]), .Z(n1971) );
  ND2 U769 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n476) );
  AN3 U770 ( .A(n224), .B(n279), .C(input_log2[45]), .Z(n1970) );
  AN3 U771 ( .A(n475), .B(n278), .C(input_log2[44]), .Z(n1969) );
  EO U772 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n475) );
  EO U773 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1102) );
  AN3 U774 ( .A(n371), .B(n279), .C(input_log2[43]), .Z(n1896) );
  NR3 U775 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n371) );
  AN3 U776 ( .A(n373), .B(n278), .C(input_log2[44]), .Z(n1895) );
  AO4 U777 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n373) );
  AN3 U778 ( .A(n370), .B(input_log2[45]), .C(input_log2[44]), .Z(n1894) );
  ND3 U779 ( .A(n224), .B(n225), .C(n223), .Z(n370) );
  AN3 U780 ( .A(n372), .B(n279), .C(input_log2[45]), .Z(n1892) );
  ND2 U781 ( .A(n223), .B(n224), .Z(n372) );
  AN3 U782 ( .A(n223), .B(n278), .C(input_log2[44]), .Z(n1904) );
  AN3 U783 ( .A(n344), .B(n277), .C(input_log2[45]), .Z(n1903) );
  NR3 U784 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n344) );
  AN3 U785 ( .A(input_log2[44]), .B(n264), .C(input_log2[43]), .Z(n2024) );
  AN3 U786 ( .A(n329), .B(input_log2[45]), .C(input_log2[43]), .Z(n2023) );
  ND3 U787 ( .A(n224), .B(n225), .C(n223), .Z(n329) );
  AN3 U788 ( .A(n332), .B(n278), .C(input_log2[43]), .Z(n2022) );
  ND3 U789 ( .A(n224), .B(n225), .C(n223), .Z(n332) );
  AN3 U790 ( .A(n331), .B(n277), .C(input_log2[44]), .Z(n2020) );
  AO4 U791 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n331) );
  AN3 U792 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .Z(
        n533) );
  EN U793 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n511) );
  EO U794 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n468) );
  EN U795 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n436) );
  EO U796 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n434) );
  EO U797 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n450) );
  EO U798 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n445) );
  EO U799 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n403) );
  EO U800 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n418) );
  EO U801 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n416) );
  EO U802 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n391) );
  EO U803 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n393) );
  EN U804 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n395) );
  EO U805 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n362) );
  EN U806 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n365) );
  EN U807 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n364) );
  ND3 U808 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n1775) );
  ND3 U809 ( .A(n278), .B(n279), .C(input_log2[43]), .Z(n2061) );
  ND3 U810 ( .A(n278), .B(n279), .C(n559), .Z(n2062) );
  AO4 U811 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[41]), .Z(n559) );
  ND3 U812 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n842) );
  ND3 U813 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n838) );
  ND3 U814 ( .A(n1392), .B(n1391), .C(n1390), .Z(n846) );
  ND2 U815 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1392) );
  ND2 U816 ( .A(input_log2[40]), .B(n223), .Z(n1391) );
  ND2 U817 ( .A(input_log2[41]), .B(n223), .Z(n1390) );
  ND3 U818 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n805) );
  ND3 U819 ( .A(n224), .B(n225), .C(input_log2[42]), .Z(n825) );
  ND3 U820 ( .A(n1474), .B(n1473), .C(n1472), .Z(n785) );
  ND2 U821 ( .A(input_log2[42]), .B(n225), .Z(n1474) );
  ND2 U822 ( .A(n224), .B(n225), .Z(n1473) );
  ND2 U823 ( .A(input_log2[42]), .B(n224), .Z(n1472) );
  ND3 U824 ( .A(input_log2[42]), .B(n224), .C(input_log2[40]), .Z(n763) );
  ND3 U825 ( .A(n2056), .B(n2055), .C(n2054), .Z(n570) );
  MUX21L U826 ( .A(n2051), .B(n2050), .S(input_log2[44]), .Z(n2056) );
  MUX21L U827 ( .A(n2048), .B(n2049), .S(input_log2[45]), .Z(n2055) );
  MUX21L U828 ( .A(n2052), .B(n2053), .S(input_log2[45]), .Z(n2054) );
  ND3 U829 ( .A(n265), .B(n279), .C(input_log2[45]), .Z(n1995) );
  ND3 U830 ( .A(n278), .B(n279), .C(n591), .Z(n1881) );
  AO7 U831 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n591) );
  ND3 U832 ( .A(n1410), .B(n1409), .C(n1408), .Z(n640) );
  ND2 U833 ( .A(input_log2[42]), .B(n225), .Z(n1410) );
  ND2 U834 ( .A(n224), .B(n225), .Z(n1409) );
  ND2 U835 ( .A(input_log2[42]), .B(n224), .Z(n1408) );
  ND3 U836 ( .A(n1461), .B(n1460), .C(n1459), .Z(n669) );
  ND2 U837 ( .A(input_log2[41]), .B(n225), .Z(n1461) );
  ND2 U838 ( .A(input_log2[42]), .B(n225), .Z(n1460) );
  ND2 U839 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1459) );
  ND3 U840 ( .A(n1224), .B(n1223), .C(n1222), .Z(n662) );
  ND2 U841 ( .A(input_log2[42]), .B(n225), .Z(n1224) );
  ND2 U842 ( .A(n224), .B(n225), .Z(n1223) );
  ND2 U843 ( .A(input_log2[42]), .B(n224), .Z(n1222) );
  ND3 U844 ( .A(n223), .B(n225), .C(input_log2[41]), .Z(n896) );
  ND3 U845 ( .A(n1573), .B(n1572), .C(n1571), .Z(n914) );
  ND2 U846 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1573) );
  ND2 U847 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1572) );
  ND2 U848 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1571) );
  ND3 U849 ( .A(input_log2[43]), .B(n308), .C(input_log2[44]), .Z(n2089) );
  ND3 U850 ( .A(n224), .B(n225), .C(n223), .Z(n308) );
  ND3 U851 ( .A(n310), .B(n278), .C(input_log2[44]), .Z(n2090) );
  ND2 U852 ( .A(n1758), .B(n1757), .Z(n310) );
  ND2 U853 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1758) );
  ND2 U854 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1757) );
  ND3 U855 ( .A(n303), .B(n277), .C(n279), .Z(n2099) );
  ND2 U856 ( .A(n1846), .B(n223), .Z(n303) );
  EO U857 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1846) );
  ND3 U858 ( .A(n1750), .B(n1749), .C(n1748), .Z(n522) );
  ND2 U859 ( .A(input_log2[41]), .B(n225), .Z(n1750) );
  ND2 U860 ( .A(input_log2[42]), .B(n225), .Z(n1749) );
  ND2 U861 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1748) );
  ND3 U862 ( .A(n1044), .B(n1043), .C(n1042), .Z(n467) );
  ND2 U863 ( .A(input_log2[40]), .B(n224), .Z(n1044) );
  ND2 U864 ( .A(n223), .B(n224), .Z(n1043) );
  ND2 U865 ( .A(input_log2[40]), .B(n223), .Z(n1042) );
  ND3 U866 ( .A(n1648), .B(n1647), .C(n1646), .Z(n489) );
  ND2 U867 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1648) );
  ND2 U868 ( .A(input_log2[40]), .B(n223), .Z(n1647) );
  ND2 U869 ( .A(input_log2[41]), .B(n223), .Z(n1646) );
  ND3 U870 ( .A(n223), .B(n225), .C(input_log2[41]), .Z(n461) );
  ND3 U871 ( .A(n1138), .B(n1137), .C(n1136), .Z(n407) );
  ND2 U872 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1138) );
  ND2 U873 ( .A(input_log2[40]), .B(n223), .Z(n1137) );
  ND2 U874 ( .A(input_log2[41]), .B(n223), .Z(n1136) );
  ND3 U875 ( .A(n1818), .B(n1817), .C(n1816), .Z(n431) );
  ND2 U876 ( .A(input_log2[41]), .B(n225), .Z(n1818) );
  ND2 U877 ( .A(n223), .B(n225), .Z(n1817) );
  ND2 U878 ( .A(input_log2[41]), .B(n223), .Z(n1816) );
  ND3 U879 ( .A(n1444), .B(n1443), .C(n1442), .Z(n387) );
  ND2 U880 ( .A(input_log2[42]), .B(n225), .Z(n1444) );
  ND2 U881 ( .A(n224), .B(n225), .Z(n1443) );
  ND2 U882 ( .A(input_log2[42]), .B(n224), .Z(n1442) );
  ND3 U883 ( .A(n1612), .B(n1611), .C(n1610), .Z(n394) );
  ND2 U884 ( .A(input_log2[41]), .B(n225), .Z(n1612) );
  ND2 U885 ( .A(n223), .B(n225), .Z(n1611) );
  ND2 U886 ( .A(input_log2[41]), .B(n223), .Z(n1610) );
  ND3 U887 ( .A(n349), .B(n277), .C(input_log2[45]), .Z(n1948) );
  AO7 U888 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n349) );
  ND3 U889 ( .A(n333), .B(n277), .C(n279), .Z(n2026) );
  NR3 U890 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n333) );
  AO4 U891 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n497) );
  AO4 U892 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n348) );
  AO7 U893 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n319) );
  NR2 U894 ( .A(input_log2[42]), .B(n224), .Z(n576) );
  ND2 U895 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1511) );
  ND2 U896 ( .A(input_log2[42]), .B(n225), .Z(n1322) );
  ND2 U897 ( .A(input_log2[40]), .B(n224), .Z(n1557) );
  ND2 U898 ( .A(input_log2[41]), .B(n223), .Z(n1779) );
  ND2 U899 ( .A(input_log2[40]), .B(n223), .Z(n1776) );
  ND2 U900 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1655) );
  ND2 U901 ( .A(input_log2[41]), .B(n223), .Z(n1537) );
  ND2 U902 ( .A(input_log2[40]), .B(n223), .Z(n1538) );
  ND2 U903 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1103) );
  ND2 U904 ( .A(input_log2[42]), .B(n224), .Z(n1439) );
  ND2 U905 ( .A(input_log2[40]), .B(n223), .Z(n1402) );
  ND2 U906 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1543) );
  ND2 U907 ( .A(n579), .B(n279), .Z(n1922) );
  AO4 U908 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n579) );
  ND2 U909 ( .A(n1745), .B(n1744), .Z(n587) );
  ND2 U910 ( .A(n223), .B(n224), .Z(n1744) );
  EO U911 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1745) );
  ND2 U912 ( .A(n1640), .B(n1639), .Z(n584) );
  MUX21L U913 ( .A(input_log2[42]), .B(n1638), .S(input_log2[40]), .Z(n1640)
         );
  ND2 U914 ( .A(input_log2[42]), .B(n224), .Z(n1639) );
  NR2 U915 ( .A(input_log2[42]), .B(n224), .Z(n1638) );
  ND2 U916 ( .A(n1807), .B(n1806), .Z(n589) );
  MUX21L U917 ( .A(n225), .B(n1805), .S(input_log2[42]), .Z(n1807) );
  ND2 U918 ( .A(input_log2[41]), .B(n223), .Z(n1806) );
  NR2 U919 ( .A(input_log2[41]), .B(n225), .Z(n1805) );
  ND2 U920 ( .A(n1631), .B(n223), .Z(n583) );
  ND2 U921 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1631) );
  ND2 U922 ( .A(n1664), .B(n1663), .Z(n585) );
  MUX21L U923 ( .A(n224), .B(n1662), .S(input_log2[42]), .Z(n1664) );
  ND2 U924 ( .A(input_log2[40]), .B(n224), .Z(n1663) );
  NR2 U925 ( .A(input_log2[40]), .B(n224), .Z(n1662) );
  ND2 U926 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1212) );
  ND2 U927 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1107) );
  ND2 U928 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1108) );
  ND2 U929 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1105) );
  ND2 U930 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1106) );
  ND2 U931 ( .A(input_log2[42]), .B(n224), .Z(n1406) );
  ND2 U932 ( .A(input_log2[42]), .B(n224), .Z(n1234) );
  ND2 U933 ( .A(input_log2[42]), .B(n224), .Z(n1049) );
  ND2 U934 ( .A(input_log2[42]), .B(n224), .Z(n1081) );
  ND2 U935 ( .A(input_log2[41]), .B(n223), .Z(n961) );
  ND2 U936 ( .A(input_log2[42]), .B(n225), .Z(n963) );
  ND2 U937 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n964) );
  ND2 U938 ( .A(input_log2[41]), .B(n225), .Z(n988) );
  ND2 U939 ( .A(input_log2[40]), .B(n224), .Z(n1799) );
  ND2 U940 ( .A(input_log2[42]), .B(n225), .Z(n1614) );
  ND2 U941 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1413) );
  ND2 U942 ( .A(input_log2[41]), .B(n223), .Z(n1414) );
  ND2 U943 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1556) );
  ND2 U944 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1465) );
  ND2 U945 ( .A(input_log2[44]), .B(n278), .Z(n2059) );
  ND2 U946 ( .A(n279), .B(n565), .Z(n2096) );
  ND2 U947 ( .A(n1810), .B(n1809), .Z(n565) );
  MUX21L U948 ( .A(n225), .B(n1808), .S(input_log2[42]), .Z(n1810) );
  ND2 U949 ( .A(input_log2[41]), .B(n225), .Z(n1809) );
  ND2 U950 ( .A(input_log2[42]), .B(n224), .Z(n1608) );
  ND2 U951 ( .A(input_log2[42]), .B(n225), .Z(n1698) );
  ND2 U952 ( .A(input_log2[42]), .B(n225), .Z(n1803) );
  ND2 U953 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1210) );
  ND2 U954 ( .A(input_log2[41]), .B(n223), .Z(n1327) );
  ND2 U955 ( .A(input_log2[41]), .B(n225), .Z(n1491) );
  ND2 U956 ( .A(n1417), .B(input_log2[40]), .Z(n1420) );
  NR2 U957 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1417) );
  ND2 U958 ( .A(input_log2[42]), .B(n224), .Z(n1382) );
  ND2 U959 ( .A(input_log2[41]), .B(n223), .Z(n1116) );
  ND2 U960 ( .A(n966), .B(n965), .Z(n828) );
  ND2 U961 ( .A(input_log2[40]), .B(n223), .Z(n966) );
  ND2 U962 ( .A(input_log2[40]), .B(n224), .Z(n965) );
  ND2 U963 ( .A(n1160), .B(n1159), .Z(n836) );
  MUX21L U964 ( .A(n225), .B(n1158), .S(input_log2[42]), .Z(n1160) );
  ND2 U965 ( .A(n224), .B(n225), .Z(n1159) );
  ND2 U966 ( .A(n1181), .B(n1180), .Z(n837) );
  MUX21L U967 ( .A(n1178), .B(n1179), .S(input_log2[40]), .Z(n1181) );
  ND2 U968 ( .A(n1177), .B(input_log2[40]), .Z(n1180) );
  ND2 U969 ( .A(input_log2[42]), .B(n224), .Z(n850) );
  ND2 U970 ( .A(n1404), .B(n1403), .Z(n847) );
  ND2 U971 ( .A(n223), .B(n224), .Z(n1404) );
  ND2 U972 ( .A(input_log2[40]), .B(n223), .Z(n1403) );
  ND2 U973 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n845) );
  ND2 U974 ( .A(n1464), .B(n225), .Z(n848) );
  EO U975 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1464) );
  ND2 U976 ( .A(n1048), .B(input_log2[42]), .Z(n865) );
  EO U977 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1048) );
  ND2 U978 ( .A(input_log2[42]), .B(n225), .Z(n866) );
  ND2 U979 ( .A(n1094), .B(n1093), .Z(n867) );
  ND2 U980 ( .A(input_log2[42]), .B(n225), .Z(n1093) );
  EO U981 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1094) );
  ND2 U982 ( .A(n1601), .B(n1600), .Z(n883) );
  MUX21L U983 ( .A(n1599), .B(input_log2[41]), .S(input_log2[40]), .Z(n1601)
         );
  ND2 U984 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1600) );
  NR2 U985 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1599) );
  ND2 U986 ( .A(n1687), .B(n1686), .Z(n886) );
  MUX21L U987 ( .A(n1684), .B(n1685), .S(input_log2[42]), .Z(n1687) );
  ND2 U988 ( .A(n1683), .B(input_log2[40]), .Z(n1686) );
  NR2 U989 ( .A(input_log2[40]), .B(n224), .Z(n1684) );
  ND2 U990 ( .A(n1170), .B(input_log2[41]), .Z(n871) );
  EN U991 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1170) );
  ND2 U992 ( .A(n1193), .B(n1192), .Z(n872) );
  MUX21L U993 ( .A(n1190), .B(n1191), .S(input_log2[41]), .Z(n1193) );
  ND2 U994 ( .A(n1189), .B(n225), .Z(n1192) );
  ND2 U995 ( .A(n1341), .B(n1340), .Z(n876) );
  MUX21L U996 ( .A(n1338), .B(n1339), .S(input_log2[40]), .Z(n1341) );
  ND2 U997 ( .A(n1337), .B(input_log2[41]), .Z(n1340) );
  ND2 U998 ( .A(n1253), .B(n1252), .Z(n874) );
  ND2 U999 ( .A(input_log2[40]), .B(n223), .Z(n1252) );
  EN U1000 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1253) );
  ND2 U1001 ( .A(n1218), .B(n1217), .Z(n873) );
  MUX21L U1002 ( .A(n1213), .B(n1214), .S(input_log2[41]), .Z(n1218) );
  MUX21L U1003 ( .A(n1215), .B(n1216), .S(input_log2[40]), .Z(n1217) );
  ND2 U1004 ( .A(n1351), .B(n1350), .Z(n877) );
  MUX21L U1005 ( .A(n1348), .B(n1349), .S(input_log2[42]), .Z(n1351) );
  ND2 U1006 ( .A(n1347), .B(input_log2[40]), .Z(n1350) );
  NR2 U1007 ( .A(input_log2[40]), .B(n224), .Z(n1348) );
  ND2 U1008 ( .A(n1287), .B(n1286), .Z(n806) );
  EN U1009 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1287) );
  EO U1010 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1286) );
  ND2 U1011 ( .A(n1355), .B(n1354), .Z(n809) );
  MUX21L U1012 ( .A(n1352), .B(n1353), .S(input_log2[41]), .Z(n1355) );
  ND3 U1013 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1354) );
  ND2 U1014 ( .A(n1298), .B(n1297), .Z(n807) );
  EN U1015 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1298) );
  EN U1016 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1297) );
  ND2 U1017 ( .A(n1206), .B(n1205), .Z(n804) );
  MUX21L U1018 ( .A(n225), .B(n1204), .S(input_log2[42]), .Z(n1206) );
  ND2 U1019 ( .A(n224), .B(n225), .Z(n1205) );
  ND2 U1020 ( .A(n1688), .B(input_log2[42]), .Z(n823) );
  EN U1021 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1688) );
  ND2 U1022 ( .A(input_log2[41]), .B(n223), .Z(n821) );
  ND2 U1023 ( .A(n1617), .B(n1616), .Z(n820) );
  MUX21L U1024 ( .A(n225), .B(n1615), .S(input_log2[42]), .Z(n1617) );
  ND2 U1025 ( .A(n224), .B(n225), .Z(n1616) );
  ND2 U1026 ( .A(n1723), .B(n1722), .Z(n824) );
  MUX21L U1027 ( .A(n1720), .B(n1721), .S(input_log2[42]), .Z(n1723) );
  ND2 U1028 ( .A(n1719), .B(input_log2[40]), .Z(n1722) );
  NR2 U1029 ( .A(input_log2[40]), .B(n224), .Z(n1720) );
  ND2 U1030 ( .A(n1369), .B(n1368), .Z(n781) );
  ND2 U1031 ( .A(n223), .B(n225), .Z(n1369) );
  ND2 U1032 ( .A(input_log2[41]), .B(n223), .Z(n1368) );
  ND2 U1033 ( .A(n1416), .B(n1415), .Z(n783) );
  ND2 U1034 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1416) );
  ND2 U1035 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1415) );
  ND2 U1036 ( .A(n1377), .B(n1376), .Z(n782) );
  ND2 U1037 ( .A(n224), .B(n225), .Z(n1377) );
  ND2 U1038 ( .A(input_log2[42]), .B(n224), .Z(n1376) );
  ND2 U1039 ( .A(n1513), .B(n223), .Z(n786) );
  ND2 U1040 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1513) );
  ND2 U1041 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n787) );
  ND2 U1042 ( .A(n1583), .B(n1582), .Z(n790) );
  MUX21L U1043 ( .A(n224), .B(n1581), .S(input_log2[42]), .Z(n1583) );
  ND2 U1044 ( .A(input_log2[40]), .B(n224), .Z(n1582) );
  NR2 U1045 ( .A(input_log2[40]), .B(n224), .Z(n1581) );
  ND2 U1046 ( .A(n1725), .B(n1724), .Z(n793) );
  ND2 U1047 ( .A(input_log2[40]), .B(n223), .Z(n1725) );
  ND2 U1048 ( .A(input_log2[40]), .B(n224), .Z(n1724) );
  ND2 U1049 ( .A(input_log2[41]), .B(n1788), .Z(n794) );
  ND2 U1050 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1788) );
  ND2 U1051 ( .A(n1041), .B(n1040), .Z(n713) );
  MUX21L U1052 ( .A(n1038), .B(n225), .S(input_log2[41]), .Z(n1040) );
  AO6 U1053 ( .A(input_log2[41]), .B(n223), .C(n1039), .Z(n1041) );
  ND2 U1054 ( .A(n995), .B(n994), .Z(n711) );
  MUX21L U1055 ( .A(n993), .B(n223), .S(input_log2[41]), .Z(n995) );
  ND2 U1056 ( .A(input_log2[41]), .B(n225), .Z(n994) );
  ND2 U1057 ( .A(n1092), .B(n1091), .Z(n715) );
  ND2 U1058 ( .A(input_log2[41]), .B(n223), .Z(n1091) );
  EO U1059 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1092) );
  ND2 U1060 ( .A(n1027), .B(n1026), .Z(n712) );
  MUX21L U1061 ( .A(n224), .B(n1025), .S(input_log2[42]), .Z(n1027) );
  ND2 U1062 ( .A(n224), .B(n225), .Z(n1026) );
  ND2 U1063 ( .A(n1115), .B(n1114), .Z(n716) );
  MUX21L U1064 ( .A(n1113), .B(n223), .S(input_log2[40]), .Z(n1115) );
  ND2 U1065 ( .A(input_log2[40]), .B(n224), .Z(n1114) );
  ND2 U1066 ( .A(input_log2[42]), .B(n1645), .Z(n732) );
  ND2 U1067 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1645) );
  ND2 U1068 ( .A(n1770), .B(n1769), .Z(n735) );
  ND2 U1069 ( .A(n223), .B(n225), .Z(n1770) );
  ND2 U1070 ( .A(input_log2[41]), .B(n223), .Z(n1769) );
  ND2 U1071 ( .A(n1830), .B(n1829), .Z(n736) );
  MUX21L U1072 ( .A(n1828), .B(input_log2[41]), .S(input_log2[40]), .Z(n1830)
         );
  ND2 U1073 ( .A(input_log2[42]), .B(input_log2[40]), .Z(n1829) );
  NR2 U1074 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1828) );
  ND2 U1075 ( .A(input_log2[42]), .B(n224), .Z(n752) );
  ND2 U1076 ( .A(n1380), .B(n1379), .Z(n751) );
  MUX21L U1077 ( .A(n1378), .B(n223), .S(input_log2[40]), .Z(n1380) );
  ND2 U1078 ( .A(input_log2[40]), .B(n224), .Z(n1379) );
  ND2 U1079 ( .A(n1055), .B(n1054), .Z(n741) );
  MUX21L U1080 ( .A(n1051), .B(input_log2[42]), .S(input_log2[40]), .Z(n1054)
         );
  NR2 U1081 ( .A(n1053), .B(n1052), .Z(n1055) );
  NR2 U1082 ( .A(input_log2[42]), .B(n224), .Z(n1051) );
  ND2 U1083 ( .A(n1097), .B(n1096), .Z(n743) );
  MUX21L U1084 ( .A(n1095), .B(n225), .S(input_log2[41]), .Z(n1097) );
  ND2 U1085 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1096) );
  NR2 U1086 ( .A(input_log2[42]), .B(n225), .Z(n1095) );
  ND2 U1087 ( .A(n1071), .B(n1070), .Z(n742) );
  ND2 U1088 ( .A(input_log2[41]), .B(n223), .Z(n1071) );
  ND2 U1089 ( .A(input_log2[41]), .B(n225), .Z(n1070) );
  ND2 U1090 ( .A(n1012), .B(n1011), .Z(n739) );
  ND2 U1091 ( .A(input_log2[42]), .B(n224), .Z(n1011) );
  EO U1092 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1012) );
  ND2 U1093 ( .A(n1676), .B(n1675), .Z(n761) );
  MUX21L U1094 ( .A(n1674), .B(input_log2[40]), .S(input_log2[42]), .Z(n1676)
         );
  ND2 U1095 ( .A(input_log2[42]), .B(n224), .Z(n1675) );
  NR2 U1096 ( .A(input_log2[40]), .B(n224), .Z(n1674) );
  ND2 U1097 ( .A(n1690), .B(n1689), .Z(n762) );
  ND2 U1098 ( .A(n223), .B(n225), .Z(n1689) );
  EN U1099 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1690) );
  ND2 U1100 ( .A(n1591), .B(n1590), .Z(n599) );
  ND2 U1101 ( .A(input_log2[40]), .B(n223), .Z(n1591) );
  ND2 U1102 ( .A(input_log2[41]), .B(n223), .Z(n1590) );
  ND2 U1103 ( .A(n1774), .B(n1773), .Z(n605) );
  ND2 U1104 ( .A(input_log2[40]), .B(n223), .Z(n1773) );
  EN U1105 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1774) );
  ND2 U1106 ( .A(input_log2[40]), .B(n223), .Z(n625) );
  ND2 U1107 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n627) );
  ND2 U1108 ( .A(n1589), .B(n1588), .Z(n622) );
  MUX21L U1109 ( .A(input_log2[40]), .B(n1587), .S(input_log2[41]), .Z(n1589)
         );
  ND2 U1110 ( .A(input_log2[42]), .B(n224), .Z(n1588) );
  NR2 U1111 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1587) );
  ND2 U1112 ( .A(input_log2[42]), .B(n224), .Z(n624) );
  ND2 U1113 ( .A(n1842), .B(n1841), .Z(n628) );
  ND2 U1114 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1841) );
  EO U1115 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1842) );
  ND2 U1116 ( .A(input_log2[44]), .B(n278), .Z(n1878) );
  ND2 U1117 ( .A(n1536), .B(n1535), .Z(n643) );
  MUX21L U1118 ( .A(n1533), .B(n1534), .S(input_log2[40]), .Z(n1536) );
  ND2 U1119 ( .A(n1532), .B(input_log2[40]), .Z(n1535) );
  ND2 U1120 ( .A(n1680), .B(n1679), .Z(n648) );
  ND2 U1121 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1680) );
  ND2 U1122 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1679) );
  ND2 U1123 ( .A(n1772), .B(n1771), .Z(n651) );
  ND2 U1124 ( .A(input_log2[40]), .B(n224), .Z(n1772) );
  ND2 U1125 ( .A(input_log2[42]), .B(n224), .Z(n1771) );
  ND2 U1126 ( .A(n1531), .B(n1530), .Z(n671) );
  MUX21L U1127 ( .A(n1527), .B(input_log2[42]), .S(input_log2[40]), .Z(n1530)
         );
  NR2 U1128 ( .A(n1529), .B(n1528), .Z(n1531) );
  NR2 U1129 ( .A(input_log2[42]), .B(n224), .Z(n1527) );
  ND2 U1130 ( .A(n1289), .B(n1288), .Z(n663) );
  ND2 U1131 ( .A(n223), .B(n225), .Z(n1288) );
  EO U1132 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1289) );
  ND2 U1133 ( .A(n1147), .B(n1146), .Z(n659) );
  ND2 U1134 ( .A(input_log2[42]), .B(n225), .Z(n1146) );
  EN U1135 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1147) );
  ND2 U1136 ( .A(n1344), .B(n1343), .Z(n665) );
  ND2 U1137 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1343) );
  EN U1138 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1344) );
  ND2 U1139 ( .A(n1832), .B(n1831), .Z(n679) );
  EN U1140 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1832) );
  EO U1141 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1831) );
  ND2 U1142 ( .A(n1602), .B(n223), .Z(n674) );
  ND2 U1143 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1602) );
  ND2 U1144 ( .A(n1696), .B(n1695), .Z(n676) );
  ND2 U1145 ( .A(input_log2[40]), .B(n223), .Z(n1695) );
  EN U1146 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1696) );
  ND2 U1147 ( .A(n1066), .B(n1065), .Z(n684) );
  ND2 U1148 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1065) );
  EO U1149 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1066) );
  ND2 U1150 ( .A(n1021), .B(n1020), .Z(n683) );
  ND2 U1151 ( .A(input_log2[42]), .B(n224), .Z(n1021) );
  ND2 U1152 ( .A(input_log2[42]), .B(n225), .Z(n1020) );
  ND2 U1153 ( .A(n1085), .B(n1084), .Z(n686) );
  MUX21L U1154 ( .A(n224), .B(n1083), .S(input_log2[42]), .Z(n1085) );
  ND2 U1155 ( .A(input_log2[40]), .B(n224), .Z(n1084) );
  NR2 U1156 ( .A(input_log2[40]), .B(n224), .Z(n1083) );
  ND2 U1157 ( .A(n971), .B(n970), .Z(n681) );
  MUX21L U1158 ( .A(n969), .B(n223), .S(input_log2[40]), .Z(n971) );
  ND2 U1159 ( .A(input_log2[41]), .B(n223), .Z(n970) );
  NR2 U1160 ( .A(input_log2[41]), .B(n223), .Z(n969) );
  ND2 U1161 ( .A(n1263), .B(n1262), .Z(n692) );
  MUX21L U1162 ( .A(n1260), .B(n1261), .S(input_log2[42]), .Z(n1263) );
  ND2 U1163 ( .A(n1259), .B(n225), .Z(n1262) );
  ND2 U1164 ( .A(n1209), .B(n1208), .Z(n690) );
  MUX21L U1165 ( .A(n1207), .B(input_log2[41]), .S(input_log2[40]), .Z(n1209)
         );
  ND2 U1166 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1208) );
  NR2 U1167 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1207) );
  ND2 U1168 ( .A(n1301), .B(n1300), .Z(n693) );
  MUX21L U1169 ( .A(n225), .B(n1299), .S(input_log2[42]), .Z(n1301) );
  ND2 U1170 ( .A(input_log2[41]), .B(n223), .Z(n1300) );
  NR2 U1171 ( .A(input_log2[41]), .B(n225), .Z(n1299) );
  ND2 U1172 ( .A(n1240), .B(n1239), .Z(n691) );
  MUX21L U1173 ( .A(n1237), .B(n1238), .S(input_log2[40]), .Z(n1240) );
  ND2 U1174 ( .A(n1236), .B(input_log2[40]), .Z(n1239) );
  ND2 U1175 ( .A(n1325), .B(n1324), .Z(n694) );
  ND2 U1176 ( .A(input_log2[40]), .B(n223), .Z(n1325) );
  ND2 U1177 ( .A(input_log2[40]), .B(n224), .Z(n1324) );
  ND2 U1178 ( .A(n1694), .B(n1693), .Z(n705) );
  MUX21L U1179 ( .A(n1691), .B(n1692), .S(input_log2[41]), .Z(n1694) );
  ND3 U1180 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1693) );
  ND2 U1181 ( .A(n1790), .B(n1789), .Z(n707) );
  ND2 U1182 ( .A(n223), .B(n225), .Z(n1789) );
  EO U1183 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1790) );
  ND2 U1184 ( .A(n1743), .B(n1742), .Z(n706) );
  MUX21L U1185 ( .A(n225), .B(n1741), .S(input_log2[42]), .Z(n1743) );
  ND2 U1186 ( .A(n224), .B(n225), .Z(n1742) );
  ND2 U1187 ( .A(n1839), .B(n1838), .Z(n708) );
  EN U1188 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1839) );
  EO U1189 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1838) );
  ND2 U1190 ( .A(n1375), .B(n223), .Z(n941) );
  EN U1191 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1375) );
  ND2 U1192 ( .A(n1500), .B(n1499), .Z(n946) );
  MUX21L U1193 ( .A(n1498), .B(input_log2[40]), .S(input_log2[42]), .Z(n1500)
         );
  ND2 U1194 ( .A(input_log2[42]), .B(n224), .Z(n1499) );
  NR2 U1195 ( .A(input_log2[40]), .B(n224), .Z(n1498) );
  ND2 U1196 ( .A(n1412), .B(input_log2[42]), .Z(n943) );
  EO U1197 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1412) );
  ND2 U1198 ( .A(n1547), .B(n1546), .Z(n947) );
  MUX21L U1199 ( .A(n1545), .B(input_log2[42]), .S(input_log2[40]), .Z(n1547)
         );
  ND2 U1200 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1546) );
  NR2 U1201 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1545) );
  ND2 U1202 ( .A(n1398), .B(n1397), .Z(n942) );
  ND2 U1203 ( .A(input_log2[42]), .B(n225), .Z(n1397) );
  EO U1204 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1398) );
  ND2 U1205 ( .A(n1447), .B(n1446), .Z(n944) );
  MUX21L U1206 ( .A(n224), .B(n1445), .S(input_log2[42]), .Z(n1447) );
  ND2 U1207 ( .A(n224), .B(n225), .Z(n1446) );
  ND2 U1208 ( .A(n1553), .B(n1552), .Z(n948) );
  MUX21L U1209 ( .A(n1550), .B(n225), .S(input_log2[41]), .Z(n1552) );
  AO6 U1210 ( .A(input_log2[41]), .B(n223), .C(n1551), .Z(n1553) );
  ND2 U1211 ( .A(n960), .B(n959), .Z(n925) );
  ND2 U1212 ( .A(n223), .B(n224), .Z(n959) );
  EN U1213 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n960) );
  ND2 U1214 ( .A(input_log2[42]), .B(n225), .Z(n930) );
  ND2 U1215 ( .A(n1008), .B(n1007), .Z(n927) );
  MUX21L U1216 ( .A(n1005), .B(n1006), .S(input_log2[40]), .Z(n1008) );
  ND2 U1217 ( .A(n1004), .B(input_log2[40]), .Z(n1007) );
  ND2 U1218 ( .A(n985), .B(n223), .Z(n926) );
  ND2 U1219 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n985) );
  ND2 U1220 ( .A(n1019), .B(n1018), .Z(n928) );
  MUX21L U1221 ( .A(n1016), .B(n1017), .S(input_log2[42]), .Z(n1019) );
  ND2 U1222 ( .A(n1015), .B(n225), .Z(n1018) );
  ND2 U1223 ( .A(n1598), .B(n1597), .Z(n950) );
  ND2 U1224 ( .A(input_log2[42]), .B(n224), .Z(n1597) );
  EO U1225 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1598) );
  ND2 U1226 ( .A(n1714), .B(n1713), .Z(n954) );
  ND2 U1227 ( .A(input_log2[42]), .B(n224), .Z(n1713) );
  EO U1228 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1714) );
  ND2 U1229 ( .A(n1658), .B(n1657), .Z(n953) );
  MUX21L U1230 ( .A(n224), .B(n1656), .S(input_log2[40]), .Z(n1658) );
  ND2 U1231 ( .A(input_log2[42]), .B(n225), .Z(n1657) );
  NR2 U1232 ( .A(input_log2[42]), .B(n224), .Z(n1656) );
  ND2 U1233 ( .A(n1827), .B(n1826), .Z(n957) );
  ND2 U1234 ( .A(n223), .B(n224), .Z(n1826) );
  EO U1235 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1827) );
  ND2 U1236 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1024) );
  ND2 U1237 ( .A(input_log2[41]), .B(n225), .Z(n1109) );
  ND2 U1238 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1110) );
  ND2 U1239 ( .A(input_log2[42]), .B(n224), .Z(n1469) );
  ND2 U1240 ( .A(n987), .B(n986), .Z(n892) );
  ND2 U1241 ( .A(input_log2[41]), .B(n223), .Z(n986) );
  EN U1242 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n987) );
  ND2 U1243 ( .A(n1400), .B(n1399), .Z(n909) );
  EN U1244 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1400) );
  EO U1245 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1399) );
  ND2 U1246 ( .A(n1431), .B(n1430), .Z(n911) );
  MUX21L U1247 ( .A(n1429), .B(n223), .S(input_log2[40]), .Z(n1431) );
  ND2 U1248 ( .A(input_log2[41]), .B(n223), .Z(n1430) );
  NR2 U1249 ( .A(input_log2[41]), .B(n223), .Z(n1429) );
  ND2 U1250 ( .A(n1156), .B(n225), .Z(n899) );
  EN U1251 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1156) );
  ND2 U1252 ( .A(n1317), .B(n1316), .Z(n905) );
  MUX21L U1253 ( .A(n1314), .B(n1315), .S(input_log2[41]), .Z(n1317) );
  ND3 U1254 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1316) );
  ND2 U1255 ( .A(input_log2[40]), .B(n1625), .Z(n917) );
  ND2 U1256 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1625) );
  ND2 U1257 ( .A(n1716), .B(n1715), .Z(n920) );
  ND2 U1258 ( .A(input_log2[42]), .B(n225), .Z(n1715) );
  EO U1259 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1716) );
  ND2 U1260 ( .A(n1673), .B(n1672), .Z(n919) );
  MUX21L U1261 ( .A(n1671), .B(input_log2[40]), .S(input_log2[42]), .Z(n1673)
         );
  ND2 U1262 ( .A(input_log2[42]), .B(n224), .Z(n1672) );
  NR2 U1263 ( .A(input_log2[40]), .B(n224), .Z(n1671) );
  ND2 U1264 ( .A(n1764), .B(n1763), .Z(n922) );
  ND2 U1265 ( .A(n224), .B(n225), .Z(n1764) );
  ND2 U1266 ( .A(input_log2[42]), .B(n225), .Z(n1763) );
  ND2 U1267 ( .A(input_log2[40]), .B(n1747), .Z(n921) );
  ND2 U1268 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1747) );
  ND2 U1269 ( .A(n1840), .B(n225), .Z(n923) );
  EO U1270 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1840) );
  ND2 U1271 ( .A(input_log2[42]), .B(n224), .Z(n1128) );
  ND2 U1272 ( .A(input_log2[40]), .B(n224), .Z(n1129) );
  ND2 U1273 ( .A(input_log2[42]), .B(n224), .Z(n1227) );
  ND2 U1274 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1139) );
  ND2 U1275 ( .A(input_log2[41]), .B(n223), .Z(n1061) );
  ND2 U1276 ( .A(n1267), .B(n225), .Z(n1270) );
  NR2 U1277 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1267) );
  ND2 U1278 ( .A(input_log2[40]), .B(n224), .Z(n1171) );
  ND2 U1279 ( .A(input_log2[41]), .B(n223), .Z(n1283) );
  ND2 U1280 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1291) );
  ND2 U1281 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1796) );
  ND2 U1282 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1682) );
  ND2 U1283 ( .A(input_log2[45]), .B(n279), .Z(n2100) );
  ND2 U1284 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1761) );
  ND2 U1285 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1762) );
  ND2 U1286 ( .A(input_log2[42]), .B(input_log2[40]), .Z(n1242) );
  ND2 U1287 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n306) );
  ND2 U1288 ( .A(input_log2[42]), .B(n224), .Z(n1078) );
  ND2 U1289 ( .A(input_log2[41]), .B(n225), .Z(n1022) );
  ND2 U1290 ( .A(input_log2[41]), .B(n223), .Z(n1023) );
  ND2 U1291 ( .A(input_log2[42]), .B(n224), .Z(n1046) );
  ND2 U1292 ( .A(input_log2[41]), .B(n223), .Z(n1002) );
  ND2 U1293 ( .A(n1386), .B(n1385), .Z(n540) );
  MUX21L U1294 ( .A(n1384), .B(n223), .S(input_log2[40]), .Z(n1386) );
  ND2 U1295 ( .A(input_log2[40]), .B(n224), .Z(n1385) );
  ND2 U1296 ( .A(n1514), .B(n223), .Z(n544) );
  EO U1297 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1514) );
  ND2 U1298 ( .A(input_log2[41]), .B(n223), .Z(n542) );
  ND2 U1299 ( .A(n1562), .B(n1561), .Z(n545) );
  MUX21L U1300 ( .A(n1559), .B(n1560), .S(input_log2[41]), .Z(n1562) );
  ND3 U1301 ( .A(input_log2[41]), .B(n223), .C(input_log2[40]), .Z(n1561) );
  ND2 U1302 ( .A(n1166), .B(n1165), .Z(n531) );
  ND2 U1303 ( .A(input_log2[42]), .B(n225), .Z(n1165) );
  EO U1304 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1166) );
  ND2 U1305 ( .A(n1363), .B(n1362), .Z(n537) );
  ND2 U1306 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1363) );
  ND2 U1307 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1362) );
  ND2 U1308 ( .A(n1185), .B(n1184), .Z(n532) );
  ND2 U1309 ( .A(n223), .B(n225), .Z(n1184) );
  EO U1310 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1185) );
  ND2 U1311 ( .A(n1266), .B(n1265), .Z(n535) );
  MUX21L U1312 ( .A(n1264), .B(n223), .S(input_log2[41]), .Z(n1266) );
  ND2 U1313 ( .A(input_log2[41]), .B(n225), .Z(n1265) );
  ND2 U1314 ( .A(n1226), .B(n1225), .Z(n534) );
  ND2 U1315 ( .A(input_log2[42]), .B(n225), .Z(n1225) );
  EN U1316 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1226) );
  ND2 U1317 ( .A(n1704), .B(n1703), .Z(n551) );
  MUX21L U1318 ( .A(n1701), .B(n225), .S(input_log2[41]), .Z(n1703) );
  AO6 U1319 ( .A(input_log2[41]), .B(n223), .C(n1702), .Z(n1704) );
  ND2 U1320 ( .A(n1837), .B(n1836), .Z(n554) );
  MUX21L U1321 ( .A(n224), .B(n1833), .S(input_log2[40]), .Z(n1836) );
  NR2 U1322 ( .A(n1835), .B(n1834), .Z(n1837) );
  ND2 U1323 ( .A(n1515), .B(n223), .Z(n513) );
  ND2 U1324 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1515) );
  ND2 U1325 ( .A(n1424), .B(n1423), .Z(n510) );
  ND2 U1326 ( .A(input_log2[42]), .B(n224), .Z(n1423) );
  EO U1327 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1424) );
  ND2 U1328 ( .A(n1619), .B(n225), .Z(n518) );
  EN U1329 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1619) );
  ND2 U1330 ( .A(input_log2[41]), .B(n225), .Z(n520) );
  ND2 U1331 ( .A(n1718), .B(n1717), .Z(n521) );
  ND2 U1332 ( .A(n223), .B(n225), .Z(n1717) );
  EO U1333 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1718) );
  ND2 U1334 ( .A(n1478), .B(n1477), .Z(n482) );
  MUX21L U1335 ( .A(n1476), .B(n223), .S(input_log2[40]), .Z(n1478) );
  ND2 U1336 ( .A(input_log2[40]), .B(n224), .Z(n1477) );
  ND2 U1337 ( .A(n1542), .B(n1541), .Z(n484) );
  MUX21L U1338 ( .A(n224), .B(n1540), .S(input_log2[42]), .Z(n1542) );
  ND2 U1339 ( .A(n224), .B(n225), .Z(n1541) );
  ND2 U1340 ( .A(n1401), .B(n223), .Z(n479) );
  ND2 U1341 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1401) );
  ND2 U1342 ( .A(n1453), .B(n1452), .Z(n481) );
  MUX21L U1343 ( .A(n224), .B(n1451), .S(input_log2[42]), .Z(n1453) );
  ND2 U1344 ( .A(n224), .B(n225), .Z(n1452) );
  ND2 U1345 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n485) );
  ND2 U1346 ( .A(n1100), .B(n1099), .Z(n469) );
  MUX21L U1347 ( .A(n1098), .B(n225), .S(input_log2[42]), .Z(n1100) );
  ND2 U1348 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1099) );
  NR2 U1349 ( .A(input_log2[41]), .B(n225), .Z(n1098) );
  ND2 U1350 ( .A(n974), .B(n973), .Z(n465) );
  MUX21L U1351 ( .A(n972), .B(n225), .S(input_log2[41]), .Z(n974) );
  ND2 U1352 ( .A(input_log2[42]), .B(n225), .Z(n973) );
  NR2 U1353 ( .A(input_log2[42]), .B(n225), .Z(n972) );
  ND2 U1354 ( .A(n1030), .B(n1029), .Z(n466) );
  MUX21L U1355 ( .A(n225), .B(n1028), .S(input_log2[42]), .Z(n1030) );
  ND2 U1356 ( .A(n224), .B(n225), .Z(n1029) );
  ND2 U1357 ( .A(n1142), .B(n1141), .Z(n470) );
  EN U1358 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1142) );
  EO U1359 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1141) );
  ND2 U1360 ( .A(n1603), .B(n223), .Z(n487) );
  ND2 U1361 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1603) );
  ND2 U1362 ( .A(n1624), .B(n1623), .Z(n488) );
  MUX21L U1363 ( .A(n1621), .B(n1622), .S(input_log2[40]), .Z(n1624) );
  ND2 U1364 ( .A(n1620), .B(input_log2[41]), .Z(n1623) );
  ND2 U1365 ( .A(n1667), .B(n1666), .Z(n490) );
  MUX21L U1366 ( .A(n1665), .B(n223), .S(input_log2[41]), .Z(n1667) );
  ND2 U1367 ( .A(input_log2[41]), .B(n225), .Z(n1666) );
  ND2 U1368 ( .A(n1783), .B(n1782), .Z(n493) );
  ND2 U1369 ( .A(input_log2[42]), .B(n224), .Z(n1782) );
  EN U1370 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1783) );
  ND2 U1371 ( .A(n1090), .B(n1089), .Z(n438) );
  MUX21L U1372 ( .A(n1087), .B(n1088), .S(input_log2[42]), .Z(n1090) );
  ND2 U1373 ( .A(n1086), .B(n225), .Z(n1089) );
  ND2 U1374 ( .A(n976), .B(n975), .Z(n433) );
  ND2 U1375 ( .A(input_log2[40]), .B(n224), .Z(n976) );
  ND2 U1376 ( .A(input_log2[42]), .B(n224), .Z(n975) );
  ND2 U1377 ( .A(n1480), .B(n1479), .Z(n452) );
  ND2 U1378 ( .A(input_log2[41]), .B(n223), .Z(n1480) );
  ND2 U1379 ( .A(input_log2[41]), .B(n225), .Z(n1479) );
  ND2 U1380 ( .A(n1549), .B(n1548), .Z(n454) );
  ND2 U1381 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1548) );
  EO U1382 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1549) );
  ND2 U1383 ( .A(n1396), .B(n1395), .Z(n449) );
  ND2 U1384 ( .A(input_log2[41]), .B(n223), .Z(n1395) );
  EO U1385 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1396) );
  ND2 U1386 ( .A(n1506), .B(n1505), .Z(n453) );
  MUX21L U1387 ( .A(n1504), .B(n223), .S(input_log2[41]), .Z(n1506) );
  ND2 U1388 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1505) );
  NR2 U1389 ( .A(input_log2[40]), .B(n223), .Z(n1504) );
  ND2 U1390 ( .A(n1463), .B(n1462), .Z(n451) );
  ND2 U1391 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1462) );
  EN U1392 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1463) );
  ND2 U1393 ( .A(n1168), .B(n1167), .Z(n441) );
  EN U1394 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1168) );
  EO U1395 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1167) );
  ND2 U1396 ( .A(n1200), .B(n1199), .Z(n443) );
  MUX21L U1397 ( .A(n1195), .B(n1196), .S(input_log2[41]), .Z(n1200) );
  MUX21L U1398 ( .A(n1197), .B(n1198), .S(input_log2[40]), .Z(n1199) );
  ND2 U1399 ( .A(n1176), .B(n1175), .Z(n442) );
  MUX21L U1400 ( .A(n1173), .B(n1174), .S(input_log2[42]), .Z(n1176) );
  ND2 U1401 ( .A(n1172), .B(n225), .Z(n1175) );
  ND2 U1402 ( .A(n1309), .B(n1308), .Z(n446) );
  MUX21L U1403 ( .A(n225), .B(n1307), .S(input_log2[42]), .Z(n1309) );
  ND2 U1404 ( .A(n224), .B(n225), .Z(n1308) );
  ND2 U1405 ( .A(n1232), .B(n1231), .Z(n444) );
  MUX21L U1406 ( .A(input_log2[40]), .B(n1229), .S(input_log2[41]), .Z(n1231)
         );
  AO6 U1407 ( .A(input_log2[40]), .B(n223), .C(n1230), .Z(n1232) );
  NR2 U1408 ( .A(input_log2[40]), .B(n223), .Z(n1229) );
  ND2 U1409 ( .A(n1332), .B(n1331), .Z(n447) );
  MUX21L U1410 ( .A(n1330), .B(n223), .S(input_log2[40]), .Z(n1332) );
  ND2 U1411 ( .A(input_log2[40]), .B(n224), .Z(n1331) );
  ND2 U1412 ( .A(n978), .B(n977), .Z(n401) );
  ND2 U1413 ( .A(input_log2[40]), .B(n223), .Z(n978) );
  ND2 U1414 ( .A(input_log2[41]), .B(n223), .Z(n977) );
  ND2 U1415 ( .A(n1482), .B(n1481), .Z(n422) );
  ND2 U1416 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1481) );
  EN U1417 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1482) );
  ND2 U1418 ( .A(n1427), .B(n1426), .Z(n420) );
  MUX21L U1419 ( .A(n1425), .B(input_log2[41]), .S(input_log2[40]), .Z(n1427)
         );
  ND2 U1420 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1426) );
  NR2 U1421 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1425) );
  ND2 U1422 ( .A(n1458), .B(n1457), .Z(n421) );
  MUX21L U1423 ( .A(n1454), .B(input_log2[42]), .S(input_log2[40]), .Z(n1457)
         );
  NR2 U1424 ( .A(n1456), .B(n1455), .Z(n1458) );
  NR2 U1425 ( .A(input_log2[42]), .B(n224), .Z(n1454) );
  ND2 U1426 ( .A(n1524), .B(n1523), .Z(n424) );
  MUX21L U1427 ( .A(n1522), .B(n225), .S(input_log2[41]), .Z(n1524) );
  ND2 U1428 ( .A(input_log2[42]), .B(n225), .Z(n1523) );
  NR2 U1429 ( .A(input_log2[42]), .B(n225), .Z(n1522) );
  ND2 U1430 ( .A(n1187), .B(n1186), .Z(n410) );
  ND2 U1431 ( .A(n223), .B(n225), .Z(n1186) );
  EO U1432 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1187) );
  ND2 U1433 ( .A(n1247), .B(n1246), .Z(n412) );
  EO U1434 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1247) );
  EO U1435 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1246) );
  ND2 U1436 ( .A(n1274), .B(n1273), .Z(n413) );
  MUX21L U1437 ( .A(n224), .B(n1272), .S(input_log2[40]), .Z(n1274) );
  ND2 U1438 ( .A(input_log2[42]), .B(n224), .Z(n1273) );
  NR2 U1439 ( .A(input_log2[42]), .B(n224), .Z(n1272) );
  ND2 U1440 ( .A(n1346), .B(n1345), .Z(n415) );
  ND2 U1441 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1345) );
  EN U1442 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1346) );
  ND2 U1443 ( .A(n1652), .B(n1651), .Z(n427) );
  ND2 U1444 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1652) );
  ND2 U1445 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1651) );
  ND2 U1446 ( .A(n1630), .B(n1629), .Z(n426) );
  MUX21L U1447 ( .A(n1626), .B(input_log2[42]), .S(input_log2[41]), .Z(n1629)
         );
  NR2 U1448 ( .A(n1628), .B(n1627), .Z(n1630) );
  NR2 U1449 ( .A(input_log2[42]), .B(n225), .Z(n1626) );
  ND2 U1450 ( .A(n1374), .B(n1373), .Z(n384) );
  MUX21L U1451 ( .A(n1372), .B(n223), .S(input_log2[40]), .Z(n1374) );
  ND2 U1452 ( .A(input_log2[41]), .B(n223), .Z(n1373) );
  NR2 U1453 ( .A(input_log2[41]), .B(n223), .Z(n1372) );
  ND2 U1454 ( .A(n1485), .B(n1484), .Z(n388) );
  MUX21L U1455 ( .A(n1483), .B(n225), .S(input_log2[41]), .Z(n1485) );
  ND2 U1456 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1484) );
  NR2 U1457 ( .A(input_log2[42]), .B(n225), .Z(n1483) );
  ND2 U1458 ( .A(n1497), .B(n1496), .Z(n389) );
  MUX21L U1459 ( .A(n224), .B(n1495), .S(input_log2[40]), .Z(n1497) );
  ND2 U1460 ( .A(input_log2[42]), .B(n224), .Z(n1496) );
  NR2 U1461 ( .A(input_log2[42]), .B(n224), .Z(n1495) );
  ND2 U1462 ( .A(n1169), .B(n223), .Z(n375) );
  ND2 U1463 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1169) );
  ND2 U1464 ( .A(n1290), .B(n223), .Z(n379) );
  ND2 U1465 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1290) );
  ND2 U1466 ( .A(n1335), .B(n1334), .Z(n381) );
  MUX21L U1467 ( .A(n1333), .B(n223), .S(input_log2[40]), .Z(n1335) );
  ND2 U1468 ( .A(input_log2[41]), .B(n223), .Z(n1334) );
  NR2 U1469 ( .A(input_log2[41]), .B(n223), .Z(n1333) );
  ND2 U1470 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n376) );
  ND2 U1471 ( .A(n1304), .B(n1303), .Z(n380) );
  ND2 U1472 ( .A(input_log2[42]), .B(n225), .Z(n1303) );
  EN U1473 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1304) );
  ND2 U1474 ( .A(n1249), .B(n1248), .Z(n378) );
  ND2 U1475 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1249) );
  ND2 U1476 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1248) );
  ND2 U1477 ( .A(n1358), .B(n1357), .Z(n382) );
  MUX21L U1478 ( .A(n1356), .B(n223), .S(input_log2[40]), .Z(n1358) );
  ND2 U1479 ( .A(input_log2[41]), .B(n223), .Z(n1357) );
  NR2 U1480 ( .A(input_log2[41]), .B(n223), .Z(n1356) );
  ND2 U1481 ( .A(n1795), .B(n1794), .Z(n398) );
  ND2 U1482 ( .A(input_log2[40]), .B(n223), .Z(n1794) );
  EO U1483 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1795) );
  ND2 U1484 ( .A(n1735), .B(n1734), .Z(n397) );
  MUX21L U1485 ( .A(n224), .B(n1733), .S(input_log2[42]), .Z(n1735) );
  ND2 U1486 ( .A(input_log2[40]), .B(n224), .Z(n1734) );
  NR2 U1487 ( .A(input_log2[40]), .B(n224), .Z(n1733) );
  ND2 U1488 ( .A(n1845), .B(n223), .Z(n399) );
  EO U1489 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1845) );
  ND2 U1490 ( .A(n1516), .B(n223), .Z(n357) );
  ND2 U1491 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1516) );
  ND2 U1492 ( .A(n1526), .B(n1525), .Z(n358) );
  ND2 U1493 ( .A(input_log2[40]), .B(n223), .Z(n1525) );
  EN U1494 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1526) );
  ND2 U1495 ( .A(n1428), .B(n223), .Z(n355) );
  ND2 U1496 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1428) );
  ND2 U1497 ( .A(n1565), .B(n1564), .Z(n359) );
  MUX21L U1498 ( .A(n1563), .B(n223), .S(input_log2[40]), .Z(n1565) );
  ND2 U1499 ( .A(input_log2[41]), .B(n223), .Z(n1564) );
  NR2 U1500 ( .A(input_log2[41]), .B(n223), .Z(n1563) );
  ND2 U1501 ( .A(n1786), .B(n1785), .Z(n367) );
  MUX21L U1502 ( .A(n1784), .B(n223), .S(input_log2[41]), .Z(n1786) );
  ND2 U1503 ( .A(input_log2[41]), .B(n225), .Z(n1785) );
  ND2 U1504 ( .A(n1596), .B(n1595), .Z(n361) );
  MUX21L U1505 ( .A(n1594), .B(n223), .S(input_log2[40]), .Z(n1596) );
  ND2 U1506 ( .A(input_log2[41]), .B(n223), .Z(n1595) );
  NR2 U1507 ( .A(input_log2[41]), .B(n223), .Z(n1594) );
  ND2 U1508 ( .A(n1740), .B(n1739), .Z(n366) );
  MUX21L U1509 ( .A(n1737), .B(n1738), .S(input_log2[42]), .Z(n1740) );
  ND2 U1510 ( .A(n1736), .B(n224), .Z(n1739) );
  ND2 U1511 ( .A(n1643), .B(n1642), .Z(n363) );
  MUX21L U1512 ( .A(n224), .B(n1641), .S(input_log2[42]), .Z(n1643) );
  ND2 U1513 ( .A(input_log2[40]), .B(n224), .Z(n1642) );
  NR2 U1514 ( .A(input_log2[40]), .B(n224), .Z(n1641) );
  ND2 U1515 ( .A(n1820), .B(n1819), .Z(n368) );
  ND2 U1516 ( .A(n223), .B(n224), .Z(n1820) );
  ND2 U1517 ( .A(input_log2[40]), .B(n224), .Z(n1819) );
  ND2 U1518 ( .A(n1712), .B(n1711), .Z(n339) );
  MUX21L U1519 ( .A(input_log2[42]), .B(n1710), .S(input_log2[40]), .Z(n1712)
         );
  ND2 U1520 ( .A(input_log2[42]), .B(n224), .Z(n1711) );
  NR2 U1521 ( .A(input_log2[42]), .B(n224), .Z(n1710) );
  ND2 U1522 ( .A(n1654), .B(n1653), .Z(n337) );
  ND2 U1523 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1654) );
  ND2 U1524 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1653) );
  ND2 U1525 ( .A(n1754), .B(n1753), .Z(n340) );
  EO U1526 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1754) );
  EO U1527 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1753) );
  ND2 U1528 ( .A(n1670), .B(n1669), .Z(n338) );
  MUX21L U1529 ( .A(input_log2[42]), .B(n1668), .S(input_log2[40]), .Z(n1670)
         );
  ND2 U1530 ( .A(input_log2[42]), .B(n224), .Z(n1669) );
  NR2 U1531 ( .A(input_log2[42]), .B(n224), .Z(n1668) );
  ND2 U1532 ( .A(n316), .B(n279), .Z(n2033) );
  NR3 U1533 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n316) );
  ND2 U1534 ( .A(n2105), .B(n2104), .Z(n298) );
  MUX21L U1535 ( .A(n2103), .B(n296), .S(input_log2[44]), .Z(n2104) );
  AO6 U1536 ( .A(input_log2[43]), .B(input_log2[44]), .C(input_log2[45]), .Z(
        n2105) );
  ND2 U1537 ( .A(n1762), .B(n1761), .Z(n296) );
  ND2 U1538 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1329) );
  MUX41 U1539 ( .D0(n555), .D1(n538), .D2(n546), .D3(n530), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N73) );
  MUX41 U1540 ( .D0(n525), .D1(n507), .D2(n516), .D3(n502), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N72) );
  ND4 U1541 ( .A(n2181), .B(n2180), .C(n2179), .D(n2178), .Z(n507) );
  MUX41 U1542 ( .D0(n495), .D1(n477), .D2(n486), .D3(n471), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N71) );
  MUX41 U1543 ( .D0(n464), .D1(n448), .D2(n455), .D3(n440), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N70) );
  MUX41 U1544 ( .D0(n432), .D1(n417), .D2(n425), .D3(n408), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N69) );
  MUX41 U1545 ( .D0(n400), .D1(n383), .D2(n392), .D3(n374), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N68) );
  MUX41 U1546 ( .D0(n369), .D1(n352), .D2(n360), .D3(n347), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N67) );
  ND4 U1547 ( .A(n1951), .B(n1950), .C(n1949), .D(n1948), .Z(n352) );
  MUX41 U1548 ( .D0(n343), .D1(n328), .D2(n334), .D3(n326), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N66) );
  ND2 U1549 ( .A(n1928), .B(n1927), .Z(n328) );
  ND2 U1550 ( .A(n1912), .B(n1911), .Z(n326) );
  MUX41 U1551 ( .D0(n324), .D1(n314), .D2(n317), .D3(n231), .A(input_log2[47]), 
        .B(input_log2[46]), .Z(N65) );
  ND4 U1552 ( .A(n2084), .B(n2083), .C(n2082), .D(n2081), .Z(n324) );
  ND4 U1553 ( .A(n2034), .B(n2033), .C(n2032), .D(n2031), .Z(n317) );
  EN U1554 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n725) );
  IVP U1555 ( .A(n561), .Z(n2214) );
  AO4 U1556 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n561) );
  IVP U1557 ( .A(n563), .Z(n2212) );
  AO7 U1558 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n563) );
  AN2P U1559 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n281) );
  MUX21L U1560 ( .A(n1448), .B(input_log2[40]), .S(input_log2[42]), .Z(n1450)
         );
  ND2 U1561 ( .A(input_log2[42]), .B(n224), .Z(n1449) );
  ND2 U1562 ( .A(input_log2[42]), .B(n224), .Z(n1502) );
  ND2 U1563 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1501) );
  OR2 U1564 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n282) );
  OR3 U1565 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n283) );
  AN3 U1566 ( .A(input_log2[42]), .B(n225), .C(input_log2[41]), .Z(n284) );
  AN3 U1567 ( .A(n223), .B(n225), .C(input_log2[41]), .Z(n285) );
  AN3 U1568 ( .A(n223), .B(n224), .C(input_log2[40]), .Z(n286) );
  AN3 U1569 ( .A(n223), .B(n225), .C(input_log2[41]), .Z(n287) );
  OR3 U1570 ( .A(input_log2[42]), .B(input_log2[40]), .C(input_log2[41]), .Z(
        n288) );
  MUX21L U1571 ( .A(n1822), .B(n1823), .S(input_log2[42]), .Z(n1825) );
  ND2 U1572 ( .A(n1821), .B(n224), .Z(n1824) );
  MUX21L U1573 ( .A(n2085), .B(n2086), .S(input_log2[43]), .Z(n2092) );
  MUX21L U1574 ( .A(n2087), .B(n2088), .S(input_log2[43]), .Z(n2091) );
  MUX21L U1575 ( .A(n2097), .B(n301), .S(input_log2[45]), .Z(n2102) );
  MUX21L U1576 ( .A(n2098), .B(n277), .S(input_log2[45]), .Z(n2101) );
  AN3 U1577 ( .A(n224), .B(n225), .C(input_log2[42]), .Z(n289) );
  AN2P U1578 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n290) );
  AN2P U1579 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n291) );
  MUX21L U1580 ( .A(n1700), .B(input_log2[41]), .S(input_log2[42]), .Z(n586)
         );
  ND2 U1581 ( .A(input_log2[41]), .B(n225), .Z(n1700) );
  MUX21L U1582 ( .A(input_log2[40]), .B(n1405), .S(input_log2[41]), .Z(n1407)
         );
  NR2 U1583 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1405) );
  MUX21L U1584 ( .A(n1233), .B(input_log2[40]), .S(input_log2[42]), .Z(n1235)
         );
  NR2 U1585 ( .A(input_log2[40]), .B(n224), .Z(n1233) );
  MUX21L U1586 ( .A(input_log2[40]), .B(n1080), .S(input_log2[41]), .Z(n1082)
         );
  NR2 U1587 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1080) );
  MUX21L U1588 ( .A(n224), .B(n1798), .S(input_log2[42]), .Z(n1800) );
  NR2 U1589 ( .A(input_log2[40]), .B(n224), .Z(n1798) );
  MUX21L U1590 ( .A(n2058), .B(n2057), .S(input_log2[43]), .Z(n2060) );
  NR2 U1591 ( .A(input_log2[45]), .B(n266), .Z(n2058) );
  NR2 U1592 ( .A(input_log2[45]), .B(n2214), .Z(n2057) );
  MUX21L U1593 ( .A(n2093), .B(n2094), .S(input_log2[44]), .Z(n2095) );
  NR2 U1594 ( .A(input_log2[43]), .B(n2212), .Z(n2094) );
  MUX21L U1595 ( .A(input_log2[41]), .B(n1779), .S(input_log2[40]), .Z(n564)
         );
  MUX21L U1596 ( .A(n2043), .B(n2042), .S(input_log2[45]), .Z(n2045) );
  AN3 U1597 ( .A(n574), .B(n279), .C(input_log2[43]), .Z(n2042) );
  NR3 U1598 ( .A(n281), .B(input_log2[43]), .C(input_log2[44]), .Z(n2043) );
  ND2 U1599 ( .A(n1655), .B(n223), .Z(n574) );
  MUX21L U1600 ( .A(n2040), .B(n2041), .S(input_log2[43]), .Z(n2046) );
  AN3 U1601 ( .A(n573), .B(input_log2[45]), .C(input_log2[44]), .Z(n2040) );
  AN3 U1602 ( .A(n576), .B(n278), .C(input_log2[44]), .Z(n2041) );
  AO4 U1603 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n573) );
  MUX21L U1604 ( .A(n2038), .B(n2039), .S(input_log2[43]), .Z(n2047) );
  AN3 U1605 ( .A(n575), .B(n279), .C(input_log2[45]), .Z(n2038) );
  NR3 U1606 ( .A(n1775), .B(input_log2[44]), .C(input_log2[45]), .Z(n2039) );
  AO7 U1607 ( .A(input_log2[40]), .B(input_log2[41]), .C(input_log2[42]), .Z(
        n575) );
  MUX21L U1608 ( .A(n224), .B(n1607), .S(input_log2[40]), .Z(n1609) );
  NR2 U1609 ( .A(input_log2[42]), .B(n224), .Z(n1607) );
  MUX21L U1610 ( .A(n224), .B(n1697), .S(input_log2[40]), .Z(n1699) );
  NR2 U1611 ( .A(input_log2[42]), .B(n224), .Z(n1697) );
  MUX21L U1612 ( .A(n1326), .B(n223), .S(input_log2[40]), .Z(n1328) );
  NR2 U1613 ( .A(input_log2[41]), .B(n223), .Z(n1326) );
  MUX21L U1614 ( .A(n1490), .B(n223), .S(input_log2[41]), .Z(n1492) );
  MUX21L U1615 ( .A(n225), .B(n1567), .S(input_log2[42]), .Z(n1569) );
  MUX21L U1616 ( .A(n1418), .B(n1419), .S(input_log2[40]), .Z(n1421) );
  NR2 U1617 ( .A(input_log2[41]), .B(n223), .Z(n1418) );
  MUX21L U1618 ( .A(n225), .B(n1296), .S(input_log2[41]), .Z(n841) );
  ND2 U1619 ( .A(input_log2[42]), .B(n225), .Z(n1296) );
  MUX21L U1620 ( .A(n224), .B(n225), .S(input_log2[42]), .Z(n843) );
  MUX21L U1621 ( .A(n1471), .B(n1470), .S(input_log2[40]), .Z(n849) );
  ND2 U1622 ( .A(input_log2[41]), .B(n223), .Z(n1471) );
  ND2 U1623 ( .A(input_log2[42]), .B(n224), .Z(n1470) );
  MUX21L U1624 ( .A(n1555), .B(n1554), .S(input_log2[42]), .Z(n852) );
  ND2 U1625 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1555) );
  ND2 U1626 ( .A(input_log2[40]), .B(n224), .Z(n1554) );
  MUX21L U1627 ( .A(n1157), .B(n223), .S(input_log2[40]), .Z(n870) );
  ND2 U1628 ( .A(n223), .B(n224), .Z(n1157) );
  MUX21L U1629 ( .A(n2014), .B(n2013), .S(input_log2[44]), .Z(n2017) );
  AN3 U1630 ( .A(n880), .B(input_log2[45]), .C(input_log2[43]), .Z(n2014) );
  AN3 U1631 ( .A(n879), .B(input_log2[45]), .C(input_log2[43]), .Z(n2013) );
  MUX21L U1632 ( .A(n1402), .B(input_log2[40]), .S(input_log2[41]), .Z(n880)
         );
  MUX21L U1633 ( .A(n2016), .B(n2015), .S(input_log2[45]), .Z(n2018) );
  NR3 U1634 ( .A(n267), .B(input_log2[43]), .C(input_log2[44]), .Z(n2016) );
  NR3 U1635 ( .A(n268), .B(input_log2[43]), .C(input_log2[44]), .Z(n2015) );
  MUX21L U1636 ( .A(n2011), .B(n2012), .S(input_log2[44]), .Z(n2019) );
  AN3 U1637 ( .A(n881), .B(n278), .C(input_log2[43]), .Z(n2011) );
  NR3 U1638 ( .A(n269), .B(input_log2[43]), .C(input_log2[45]), .Z(n2012) );
  ND2 U1639 ( .A(input_log2[40]), .B(n1543), .Z(n881) );
  MUX21L U1640 ( .A(n225), .B(n1144), .S(input_log2[41]), .Z(n802) );
  ND2 U1641 ( .A(n223), .B(n225), .Z(n1144) );
  MUX21L U1642 ( .A(n1318), .B(input_log2[40]), .S(input_log2[42]), .Z(n808)
         );
  ND2 U1643 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1318) );
  MUX21L U1644 ( .A(n1660), .B(n1659), .S(input_log2[41]), .Z(n822) );
  ND2 U1645 ( .A(input_log2[40]), .B(n223), .Z(n1660) );
  ND2 U1646 ( .A(input_log2[42]), .B(n225), .Z(n1659) );
  MUX21L U1647 ( .A(n2112), .B(n2113), .S(input_log2[45]), .Z(n2114) );
  AN3 U1648 ( .A(n771), .B(n279), .C(input_log2[43]), .Z(n2112) );
  EN U1649 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n771) );
  MUX21L U1650 ( .A(n1433), .B(n1432), .S(input_log2[42]), .Z(n784) );
  ND2 U1651 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1433) );
  ND2 U1652 ( .A(input_log2[40]), .B(n224), .Z(n1432) );
  MUX21L U1653 ( .A(n1644), .B(n225), .S(input_log2[41]), .Z(n791) );
  ND2 U1654 ( .A(input_log2[42]), .B(n225), .Z(n1644) );
  MUX21L U1655 ( .A(input_log2[40]), .B(input_log2[41]), .S(input_log2[42]), 
        .Z(n792) );
  MUX21L U1656 ( .A(n2188), .B(n2189), .S(input_log2[45]), .Z(n2190) );
  AN3 U1657 ( .A(n728), .B(n279), .C(input_log2[43]), .Z(n2188) );
  MUX21L U1658 ( .A(input_log2[42]), .B(input_log2[40]), .S(input_log2[41]), 
        .Z(n728) );
  MUX21L U1659 ( .A(n225), .B(n968), .S(input_log2[41]), .Z(n710) );
  ND2 U1660 ( .A(n223), .B(n225), .Z(n968) );
  MUX21L U1661 ( .A(input_log2[42]), .B(n1072), .S(input_log2[40]), .Z(n714)
         );
  ND2 U1662 ( .A(input_log2[42]), .B(n224), .Z(n1072) );
  MUX21L U1663 ( .A(n1606), .B(n1605), .S(input_log2[41]), .Z(n731) );
  ND2 U1664 ( .A(n223), .B(n225), .Z(n1606) );
  ND2 U1665 ( .A(input_log2[42]), .B(n225), .Z(n1605) );
  MUX21L U1666 ( .A(input_log2[41]), .B(input_log2[42]), .S(input_log2[40]), 
        .Z(n734) );
  MUX21L U1667 ( .A(n225), .B(n967), .S(input_log2[42]), .Z(n738) );
  ND2 U1668 ( .A(input_log2[41]), .B(n225), .Z(n967) );
  MUX21L U1669 ( .A(n1112), .B(input_log2[41]), .S(input_log2[42]), .Z(n744)
         );
  ND2 U1670 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1112) );
  MUX21L U1671 ( .A(input_log2[42]), .B(n1604), .S(input_log2[40]), .Z(n759)
         );
  ND2 U1672 ( .A(input_log2[42]), .B(n224), .Z(n1604) );
  MUX21L U1673 ( .A(n1650), .B(n223), .S(input_log2[41]), .Z(n760) );
  ND2 U1674 ( .A(input_log2[40]), .B(n223), .Z(n1650) );
  MUX21L U1675 ( .A(n1802), .B(n1801), .S(input_log2[41]), .Z(n765) );
  ND2 U1676 ( .A(n223), .B(n225), .Z(n1802) );
  ND2 U1677 ( .A(input_log2[42]), .B(n225), .Z(n1801) );
  MUX21L U1678 ( .A(n1963), .B(n1962), .S(input_log2[45]), .Z(n1965) );
  NR2 U1679 ( .A(input_log2[43]), .B(n282), .Z(n1963) );
  ND2 U1680 ( .A(n1212), .B(n223), .Z(n593) );
  MUX21L U1681 ( .A(n1876), .B(n1877), .S(input_log2[45]), .Z(n1879) );
  AN3 U1682 ( .A(n279), .B(n277), .C(n223), .Z(n1877) );
  ND2 U1683 ( .A(n1108), .B(n1107), .Z(n608) );
  MUX21L U1684 ( .A(n1586), .B(input_log2[40]), .S(input_log2[42]), .Z(n646)
         );
  ND2 U1685 ( .A(input_log2[40]), .B(n224), .Z(n1586) );
  MUX21L U1686 ( .A(n1727), .B(n1726), .S(input_log2[42]), .Z(n650) );
  ND2 U1687 ( .A(input_log2[41]), .B(n225), .Z(n1727) );
  ND2 U1688 ( .A(n224), .B(n225), .Z(n1726) );
  MUX21L U1689 ( .A(n1868), .B(n1867), .S(input_log2[45]), .Z(n1873) );
  NR2 U1690 ( .A(input_log2[43]), .B(n2211), .Z(n1868) );
  NR2 U1691 ( .A(input_log2[44]), .B(n223), .Z(n1867) );
  IVP U1692 ( .A(n631), .Z(n2211) );
  MUX21L U1693 ( .A(n1871), .B(n1872), .S(input_log2[43]), .Z(n1874) );
  NR2 U1694 ( .A(input_log2[45]), .B(n279), .Z(n1871) );
  NR2 U1695 ( .A(input_log2[44]), .B(n278), .Z(n1872) );
  MUX21L U1696 ( .A(n1869), .B(n1870), .S(input_log2[44]), .Z(n1875) );
  NR2 U1697 ( .A(input_log2[43]), .B(n283), .Z(n1870) );
  ND2 U1698 ( .A(n1106), .B(n1105), .Z(n630) );
  MUX21L U1699 ( .A(n224), .B(n1302), .S(input_log2[42]), .Z(n664) );
  ND2 U1700 ( .A(n224), .B(n225), .Z(n1302) );
  MUX21L U1701 ( .A(n1194), .B(input_log2[41]), .S(input_log2[42]), .Z(n661)
         );
  ND2 U1702 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1194) );
  MUX21L U1703 ( .A(n1678), .B(n1677), .S(input_log2[40]), .Z(n675) );
  ND2 U1704 ( .A(input_log2[41]), .B(n223), .Z(n1678) );
  ND2 U1705 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1677) );
  MUX21L U1706 ( .A(n223), .B(input_log2[41]), .S(input_log2[40]), .Z(n678) );
  MUX21L U1707 ( .A(n2201), .B(n2200), .S(input_log2[44]), .Z(n2202) );
  AN3 U1708 ( .A(input_log2[45]), .B(n697), .C(input_log2[43]), .Z(n2201) );
  ND2 U1709 ( .A(n1407), .B(n1406), .Z(n697) );
  MUX21L U1710 ( .A(n1585), .B(n1584), .S(input_log2[40]), .Z(n702) );
  ND2 U1711 ( .A(n223), .B(n224), .Z(n1585) );
  ND2 U1712 ( .A(input_log2[41]), .B(n223), .Z(n1584) );
  MUX21L U1713 ( .A(input_log2[42]), .B(n1618), .S(input_log2[41]), .Z(n703)
         );
  ND2 U1714 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1618) );
  MUX21L U1715 ( .A(n225), .B(n1661), .S(input_log2[42]), .Z(n704) );
  ND2 U1716 ( .A(input_log2[41]), .B(n225), .Z(n1661) );
  MUX21L U1717 ( .A(n1468), .B(n1467), .S(input_log2[41]), .Z(n945) );
  ND2 U1718 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1468) );
  ND2 U1719 ( .A(input_log2[42]), .B(n225), .Z(n1467) );
  MUX21L U1720 ( .A(n1032), .B(n1031), .S(input_log2[41]), .Z(n929) );
  ND2 U1721 ( .A(n223), .B(n225), .Z(n1032) );
  ND2 U1722 ( .A(input_log2[42]), .B(n225), .Z(n1031) );
  MUX21L U1723 ( .A(input_log2[40]), .B(input_log2[41]), .S(input_log2[42]), 
        .Z(n932) );
  MUX21L U1724 ( .A(n1613), .B(n224), .S(input_log2[40]), .Z(n951) );
  ND2 U1725 ( .A(n223), .B(n224), .Z(n1613) );
  MUX21L U1726 ( .A(n1633), .B(n1632), .S(input_log2[42]), .Z(n952) );
  ND2 U1727 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1633) );
  ND2 U1728 ( .A(input_log2[41]), .B(n225), .Z(n1632) );
  MUX21L U1729 ( .A(n1791), .B(n223), .S(input_log2[41]), .Z(n956) );
  ND2 U1730 ( .A(n223), .B(n225), .Z(n1791) );
  MUX21L U1731 ( .A(n224), .B(input_log2[42]), .S(input_log2[40]), .Z(n900) );
  MUX21L U1732 ( .A(n1251), .B(n1250), .S(input_log2[41]), .Z(n903) );
  ND2 U1733 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1251) );
  ND2 U1734 ( .A(input_log2[42]), .B(n225), .Z(n1250) );
  MUX21L U1735 ( .A(n224), .B(input_log2[42]), .S(input_log2[40]), .Z(n916) );
  MUX21L U1736 ( .A(n223), .B(input_log2[40]), .S(input_log2[41]), .Z(n918) );
  MUX21L U1737 ( .A(n1124), .B(n1125), .S(input_log2[41]), .Z(n1126) );
  NR2 U1738 ( .A(input_log2[42]), .B(n225), .Z(n1124) );
  NR2 U1739 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1125) );
  MUX21L U1740 ( .A(n1268), .B(n1269), .S(input_log2[42]), .Z(n1271) );
  NR2 U1741 ( .A(input_log2[40]), .B(n224), .Z(n1269) );
  MUX21L U1742 ( .A(n1241), .B(input_log2[41]), .S(input_log2[40]), .Z(n1243)
         );
  NR2 U1743 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1241) );
  MUX21L U1744 ( .A(input_log2[40]), .B(n1077), .S(input_log2[41]), .Z(n1079)
         );
  NR2 U1745 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1077) );
  MUX21L U1746 ( .A(n1131), .B(input_log2[42]), .S(input_log2[40]), .Z(n1134)
         );
  NR2 U1747 ( .A(input_log2[42]), .B(n224), .Z(n1131) );
  MUX21L U1748 ( .A(input_log2[42]), .B(n1045), .S(input_log2[40]), .Z(n1047)
         );
  NR2 U1749 ( .A(input_log2[42]), .B(n224), .Z(n1045) );
  MUX21L U1750 ( .A(n1001), .B(n223), .S(input_log2[40]), .Z(n1003) );
  NR2 U1751 ( .A(input_log2[41]), .B(n223), .Z(n1001) );
  MUX21L U1752 ( .A(n1371), .B(n1370), .S(input_log2[41]), .Z(n539) );
  ND2 U1753 ( .A(input_log2[40]), .B(n223), .Z(n1371) );
  ND2 U1754 ( .A(n223), .B(n225), .Z(n1370) );
  MUX21L U1755 ( .A(n224), .B(n1475), .S(input_log2[40]), .Z(n543) );
  ND2 U1756 ( .A(input_log2[42]), .B(n224), .Z(n1475) );
  MUX21L U1757 ( .A(n1422), .B(n225), .S(input_log2[41]), .Z(n541) );
  ND2 U1758 ( .A(input_log2[42]), .B(n225), .Z(n1422) );
  MUX21L U1759 ( .A(n1342), .B(n223), .S(input_log2[40]), .Z(n536) );
  ND2 U1760 ( .A(input_log2[41]), .B(n223), .Z(n1342) );
  MUX21L U1761 ( .A(n224), .B(n1732), .S(input_log2[42]), .Z(n552) );
  ND2 U1762 ( .A(input_log2[40]), .B(n224), .Z(n1732) );
  MUX21L U1763 ( .A(n225), .B(input_log2[41]), .S(input_log2[42]), .Z(n550) );
  MUX21L U1764 ( .A(n1781), .B(n1780), .S(input_log2[42]), .Z(n553) );
  ND2 U1765 ( .A(input_log2[41]), .B(n225), .Z(n1781) );
  ND2 U1766 ( .A(n224), .B(n225), .Z(n1780) );
  MUX21L U1767 ( .A(n2124), .B(n2125), .S(input_log2[45]), .Z(n2126) );
  AN3 U1768 ( .A(n501), .B(n279), .C(input_log2[43]), .Z(n2124) );
  EN U1769 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n501) );
  MUX21L U1770 ( .A(n2177), .B(n2176), .S(input_log2[45]), .Z(n2178) );
  AN3 U1771 ( .A(input_log2[44]), .B(n506), .C(input_log2[43]), .Z(n2177) );
  AN3 U1772 ( .A(input_log2[43]), .B(input_log2[44]), .C(n503), .Z(n2176) );
  ND2 U1773 ( .A(n1271), .B(n1270), .Z(n506) );
  MUX21L U1774 ( .A(n2175), .B(n2174), .S(input_log2[45]), .Z(n2180) );
  AN3 U1775 ( .A(input_log2[40]), .B(n279), .C(input_log2[43]), .Z(n2174) );
  NR2 U1776 ( .A(input_log2[44]), .B(n270), .Z(n2175) );
  MUX21L U1777 ( .A(n2173), .B(n2172), .S(input_log2[45]), .Z(n2181) );
  AN3 U1778 ( .A(n504), .B(n277), .C(input_log2[44]), .Z(n2172) );
  NR2 U1779 ( .A(input_log2[43]), .B(input_log2[41]), .Z(n2173) );
  MUX21L U1780 ( .A(n1171), .B(input_log2[40]), .S(input_log2[42]), .Z(n504)
         );
  MUX21L U1781 ( .A(input_log2[41]), .B(n1387), .S(input_log2[40]), .Z(n509)
         );
  ND2 U1782 ( .A(input_log2[41]), .B(n223), .Z(n1387) );
  MUX21L U1783 ( .A(n223), .B(n225), .S(input_log2[41]), .Z(n512) );
  MUX21L U1784 ( .A(n225), .B(n224), .S(input_log2[42]), .Z(n514) );
  MUX21L U1785 ( .A(n1593), .B(n1592), .S(input_log2[40]), .Z(n517) );
  ND2 U1786 ( .A(n223), .B(n224), .Z(n1593) );
  ND2 U1787 ( .A(input_log2[41]), .B(n223), .Z(n1592) );
  MUX21L U1788 ( .A(n224), .B(input_log2[42]), .S(input_log2[40]), .Z(n519) );
  MUX21L U1789 ( .A(n225), .B(input_log2[42]), .S(input_log2[41]), .Z(n523) );
  MUX21L U1790 ( .A(n1493), .B(input_log2[40]), .S(input_log2[42]), .Z(n483)
         );
  ND2 U1791 ( .A(input_log2[40]), .B(n224), .Z(n1493) );
  MUX21L U1792 ( .A(n1706), .B(n1705), .S(input_log2[42]), .Z(n491) );
  ND2 U1793 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1706) );
  ND2 U1794 ( .A(input_log2[40]), .B(n224), .Z(n1705) );
  MUX21L U1795 ( .A(input_log2[42]), .B(n224), .S(input_log2[40]), .Z(n457) );
  MUX21L U1796 ( .A(n225), .B(n1707), .S(input_log2[42]), .Z(n460) );
  ND2 U1797 ( .A(n224), .B(n225), .Z(n1707) );
  MUX21L U1798 ( .A(n1649), .B(n223), .S(input_log2[40]), .Z(n458) );
  ND2 U1799 ( .A(input_log2[41]), .B(n223), .Z(n1649) );
  MUX21L U1800 ( .A(n225), .B(n224), .S(input_log2[42]), .Z(n462) );
  MUX21L U1801 ( .A(n224), .B(n1388), .S(input_log2[40]), .Z(n419) );
  ND2 U1802 ( .A(input_log2[42]), .B(n224), .Z(n1388) );
  MUX21L U1803 ( .A(n225), .B(n1494), .S(input_log2[42]), .Z(n423) );
  ND2 U1804 ( .A(input_log2[41]), .B(n225), .Z(n1494) );
  MUX21L U1805 ( .A(n1155), .B(input_log2[41]), .S(input_log2[42]), .Z(n409)
         );
  ND2 U1806 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1155) );
  MUX21L U1807 ( .A(n1202), .B(n1201), .S(input_log2[42]), .Z(n411) );
  ND2 U1808 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1202) );
  ND2 U1809 ( .A(n224), .B(n225), .Z(n1201) );
  MUX21L U1810 ( .A(n1709), .B(n1708), .S(input_log2[41]), .Z(n428) );
  ND2 U1811 ( .A(input_log2[40]), .B(n223), .Z(n1709) );
  ND2 U1812 ( .A(n223), .B(n225), .Z(n1708) );
  MUX21L U1813 ( .A(input_log2[41]), .B(input_log2[40]), .S(input_log2[42]), 
        .Z(n429) );
  MUX21L U1814 ( .A(n224), .B(n1389), .S(input_log2[42]), .Z(n385) );
  ND2 U1815 ( .A(n224), .B(n225), .Z(n1389) );
  MUX21L U1816 ( .A(n1411), .B(input_log2[41]), .S(input_log2[42]), .Z(n386)
         );
  ND2 U1817 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1411) );
  MUX21L U1818 ( .A(n1946), .B(n1947), .S(input_log2[45]), .Z(n1949) );
  AN3 U1819 ( .A(n350), .B(input_log2[44]), .C(input_log2[43]), .Z(n1946) );
  NR2 U1820 ( .A(input_log2[43]), .B(n279), .Z(n1947) );
  ND2 U1821 ( .A(n1291), .B(n223), .Z(n350) );
  MUX21L U1822 ( .A(n1944), .B(n1945), .S(input_log2[44]), .Z(n1950) );
  AN3 U1823 ( .A(n351), .B(n278), .C(input_log2[43]), .Z(n1944) );
  ND3 U1824 ( .A(n224), .B(n225), .C(n223), .Z(n351) );
  MUX21L U1825 ( .A(n1942), .B(n1943), .S(input_log2[44]), .Z(n1951) );
  NR2 U1826 ( .A(input_log2[43]), .B(n271), .Z(n1943) );
  NR3 U1827 ( .A(input_log2[43]), .B(n288), .C(input_log2[45]), .Z(n1942) );
  MUX21L U1828 ( .A(n1486), .B(n223), .S(input_log2[41]), .Z(n356) );
  ND2 U1829 ( .A(n223), .B(n225), .Z(n1486) );
  MUX21L U1830 ( .A(input_log2[42]), .B(n1787), .S(input_log2[40]), .Z(n341)
         );
  ND2 U1831 ( .A(input_log2[42]), .B(n224), .Z(n1787) );
  MUX21L U1832 ( .A(input_log2[42]), .B(input_log2[40]), .S(input_log2[41]), 
        .Z(n342) );
  MUX21L U1833 ( .A(n1908), .B(n278), .S(input_log2[44]), .Z(n1911) );
  AN3 U1834 ( .A(n325), .B(n277), .C(input_log2[45]), .Z(n1908) );
  NR2 U1835 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n325) );
  MUX21L U1836 ( .A(n1924), .B(n279), .S(input_log2[45]), .Z(n1927) );
  AN3 U1837 ( .A(input_log2[43]), .B(n327), .C(input_log2[44]), .Z(n1924) );
  ND2 U1838 ( .A(n1292), .B(n223), .Z(n327) );
  ND2 U1839 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1292) );
  MUX21L U1840 ( .A(n2030), .B(n277), .S(input_log2[45]), .Z(n2031) );
  AN3 U1841 ( .A(input_log2[44]), .B(n272), .C(input_log2[43]), .Z(n2030) );
  MUX21L U1842 ( .A(n2080), .B(n2079), .S(input_log2[44]), .Z(n2082) );
  AN3 U1843 ( .A(n321), .B(n278), .C(input_log2[43]), .Z(n2079) );
  NR3 U1844 ( .A(input_log2[45]), .B(input_log2[43]), .C(n273), .Z(n2080) );
  AO4 U1845 ( .A(input_log2[41]), .B(input_log2[42]), .C(input_log2[40]), .D(
        input_log2[42]), .Z(n321) );
  MUX21L U1846 ( .A(n2077), .B(n2078), .S(input_log2[44]), .Z(n2083) );
  AN3 U1847 ( .A(n323), .B(n278), .C(input_log2[43]), .Z(n2077) );
  AN3 U1848 ( .A(n318), .B(input_log2[43]), .C(input_log2[45]), .Z(n2078) );
  ND2 U1849 ( .A(n1797), .B(n1796), .Z(n323) );
  MUX21L U1850 ( .A(n2075), .B(n2076), .S(input_log2[43]), .Z(n2084) );
  AN3 U1851 ( .A(n320), .B(n279), .C(input_log2[45]), .Z(n2075) );
  AN3 U1852 ( .A(n319), .B(n279), .C(input_log2[45]), .Z(n2076) );
  ND2 U1853 ( .A(n1682), .B(n223), .Z(n320) );
  ND2 U1854 ( .A(n1014), .B(n1013), .Z(n768) );
  ND2 U1855 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1013) );
  EO U1856 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1014) );
  ND2 U1857 ( .A(n1150), .B(n1149), .Z(n503) );
  MUX21L U1858 ( .A(n224), .B(n1148), .S(input_log2[42]), .Z(n1150) );
  ND2 U1859 ( .A(input_log2[40]), .B(n223), .Z(n1149) );
  NR2 U1860 ( .A(input_log2[40]), .B(n224), .Z(n1148) );
  ND2 U1861 ( .A(n2133), .B(n2132), .Z(N64) );
  MUX21L U1862 ( .A(n2131), .B(n305), .S(input_log2[47]), .Z(n2132) );
  AO2 U1863 ( .A(input_log2[46]), .B(n307), .C(input_log2[46]), .D(
        input_log2[47]), .Z(n2133) );
  NR2 U1864 ( .A(input_log2[46]), .B(n274), .Z(n2131) );
  ND2 U1865 ( .A(n2037), .B(n2036), .Z(N63) );
  MUX21L U1866 ( .A(n2035), .B(input_log2[47]), .S(input_log2[46]), .Z(n2037)
         );
  ND2 U1867 ( .A(n300), .B(input_log2[47]), .Z(n2036) );
  NR2 U1868 ( .A(input_log2[47]), .B(n275), .Z(n2035) );
  ND2 U1869 ( .A(n1921), .B(n1920), .Z(N62) );
  MUX21L U1870 ( .A(n1919), .B(n220), .S(input_log2[46]), .Z(n1921) );
  ND2 U1871 ( .A(n298), .B(n220), .Z(n1920) );
  MUX21L U1872 ( .A(n224), .B(n1364), .S(input_log2[40]), .Z(n879) );
  ND2 U1873 ( .A(input_log2[42]), .B(n224), .Z(n1364) );
  MUX81P U1874 ( .D0(n342), .D1(n338), .D2(n340), .D3(n336), .D4(n341), .D5(
        n337), .D6(n339), .D7(n335), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n343) );
  MUX81P U1875 ( .D0(n359), .D1(n223), .D2(n357), .D3(n354), .D4(n358), .D5(
        n355), .D6(n356), .D7(n353), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n360) );
  MUX81P U1876 ( .D0(n368), .D1(n364), .D2(n366), .D3(n362), .D4(n367), .D5(
        n363), .D6(n365), .D7(n361), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n369) );
  MUX81P U1877 ( .D0(n382), .D1(n378), .D2(n380), .D3(n376), .D4(n381), .D5(
        n377), .D6(n379), .D7(n375), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n383) );
  MUX81P U1878 ( .D0(n391), .D1(n387), .D2(n389), .D3(n385), .D4(n390), .D5(
        n386), .D6(n388), .D7(n384), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n392) );
  MUX81P U1879 ( .D0(n399), .D1(input_log2[40]), .D2(n397), .D3(n394), .D4(
        n398), .D5(n395), .D6(n396), .D7(n393), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n400) );
  MUX81P U1880 ( .D0(n407), .D1(n403), .D2(n405), .D3(n401), .D4(n406), .D5(
        n402), .D6(n404), .D7(n223), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n408) );
  MUX81P U1881 ( .D0(n416), .D1(n412), .D2(n414), .D3(n410), .D4(n415), .D5(
        n411), .D6(n413), .D7(n409), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n417) );
  MUX81P U1882 ( .D0(input_log2[40]), .D1(n421), .D2(n423), .D3(n419), .D4(
        n424), .D5(n420), .D6(n422), .D7(n418), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n425) );
  MUX81P U1883 ( .D0(n431), .D1(n291), .D2(n429), .D3(n426), .D4(n430), .D5(
        n427), .D6(n428), .D7(input_log2[40]), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n432) );
  MUX81P U1884 ( .D0(n439), .D1(n435), .D2(n437), .D3(n433), .D4(n438), .D5(
        n434), .D6(n436), .D7(n224), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n440) );
  MUX81P U1885 ( .D0(input_log2[40]), .D1(n444), .D2(n446), .D3(n442), .D4(
        n447), .D5(n443), .D6(n445), .D7(n441), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n448) );
  MUX81P U1886 ( .D0(n290), .D1(n451), .D2(n453), .D3(n449), .D4(n454), .D5(
        n450), .D6(n452), .D7(input_log2[40]), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n455) );
  MUX81P U1887 ( .D0(n463), .D1(n459), .D2(n461), .D3(n457), .D4(n462), .D5(
        n458), .D6(n460), .D7(n456), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n464) );
  MUX81P U1888 ( .D0(n470), .D1(n466), .D2(n468), .D3(n465), .D4(n469), .D5(
        input_log2[40]), .D6(n467), .D7(n225), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n471) );
  MUX81P U1889 ( .D0(n485), .D1(n481), .D2(n483), .D3(n479), .D4(n484), .D5(
        n480), .D6(n482), .D7(n478), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n486) );
  MUX81P U1890 ( .D0(n494), .D1(n490), .D2(n492), .D3(n488), .D4(n493), .D5(
        n489), .D6(n491), .D7(n487), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n495) );
  MUX81P U1891 ( .D0(n515), .D1(n511), .D2(n513), .D3(n509), .D4(n514), .D5(
        n510), .D6(n512), .D7(n508), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n516) );
  MUX81P U1892 ( .D0(n524), .D1(n520), .D2(n522), .D3(n518), .D4(n523), .D5(
        n519), .D6(n521), .D7(n517), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n525) );
  MUX81P U1893 ( .D0(n537), .D1(n534), .D2(input_log2[40]), .D3(n532), .D4(
        n536), .D5(n533), .D6(n535), .D7(n531), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n538) );
  MUX81P U1894 ( .D0(n545), .D1(n542), .D2(n544), .D3(n540), .D4(n289), .D5(
        n541), .D6(n543), .D7(n539), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n546) );
  MUX81P U1895 ( .D0(n554), .D1(n550), .D2(n552), .D3(n548), .D4(n553), .D5(
        n549), .D6(n551), .D7(n547), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n555) );
  MUX81P U1896 ( .D0(n589), .D1(n585), .D2(n587), .D3(n583), .D4(n588), .D5(
        n584), .D6(n586), .D7(n582), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n590) );
  MUX81P U1897 ( .D0(n606), .D1(n602), .D2(n604), .D3(n600), .D4(n605), .D5(
        n601), .D6(n603), .D7(n599), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n607) );
  MUX81P U1898 ( .D0(n628), .D1(n624), .D2(n626), .D3(n623), .D4(n627), .D5(
        input_log2[40]), .D6(n625), .D7(n622), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n629) );
  MUX81P U1899 ( .D0(n223), .D1(n223), .D2(n636), .D3(n634), .D4(n637), .D5(
        n635), .D6(n232), .D7(n633), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n638) );
  MUX81P U1900 ( .D0(n644), .D1(input_log2[41]), .D2(n642), .D3(n639), .D4(
        n643), .D5(n640), .D6(n641), .D7(n223), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n645) );
  MUX81P U1901 ( .D0(n652), .D1(n648), .D2(n650), .D3(input_log2[41]), .D4(
        n651), .D5(n647), .D6(n649), .D7(n646), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n653) );
  MUX81P U1902 ( .D0(n224), .D1(n662), .D2(n664), .D3(n660), .D4(n665), .D5(
        n661), .D6(n663), .D7(n659), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n666) );
  MUX81P U1903 ( .D0(n672), .D1(n669), .D2(n670), .D3(n667), .D4(n671), .D5(
        n668), .D6(input_log2[40]), .D7(n224), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n673) );
  MUX81P U1904 ( .D0(n679), .D1(n675), .D2(n677), .D3(input_log2[40]), .D4(
        n678), .D5(n286), .D6(n676), .D7(n674), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n680) );
  MUX81P U1905 ( .D0(n687), .D1(n683), .D2(n685), .D3(n681), .D4(n686), .D5(
        n682), .D6(n684), .D7(n223), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n688) );
  MUX81P U1906 ( .D0(n225), .D1(n691), .D2(n693), .D3(input_log2[41]), .D4(
        n694), .D5(n690), .D6(n692), .D7(n689), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n695) );
  MUX81P U1907 ( .D0(n708), .D1(n704), .D2(n706), .D3(n703), .D4(n707), .D5(
        n287), .D6(n705), .D7(n702), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n709) );
  MUX81P U1908 ( .D0(n716), .D1(n712), .D2(n714), .D3(n710), .D4(n715), .D5(
        n711), .D6(n713), .D7(n224), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n717) );
  MUX81P U1909 ( .D0(n736), .D1(n733), .D2(n285), .D3(n731), .D4(n735), .D5(
        n732), .D6(n734), .D7(n730), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n737) );
  MUX81P U1910 ( .D0(n744), .D1(n740), .D2(n742), .D3(n738), .D4(n743), .D5(
        n739), .D6(n741), .D7(n225), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n745) );
  MUX81P U1911 ( .D0(n756), .D1(n753), .D2(n754), .D3(n751), .D4(n755), .D5(
        n752), .D6(n233), .D7(n750), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n757) );
  MUX81P U1912 ( .D0(n765), .D1(n761), .D2(n763), .D3(n759), .D4(n764), .D5(
        n760), .D6(n762), .D7(n758), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n766) );
  MUX81P U1913 ( .D0(n788), .D1(n784), .D2(n786), .D3(n782), .D4(n787), .D5(
        n783), .D6(n785), .D7(n781), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n789) );
  MUX81P U1914 ( .D0(n224), .D1(n792), .D2(n793), .D3(input_log2[41]), .D4(
        n794), .D5(n791), .D6(input_log2[42]), .D7(n790), .A(input_log2[45]), 
        .B(input_log2[44]), .C(input_log2[43]), .Z(n795) );
  MUX81P U1915 ( .D0(n809), .D1(n805), .D2(n807), .D3(n803), .D4(n808), .D5(
        n804), .D6(n806), .D7(n802), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n810) );
  MUX81P U1916 ( .D0(n817), .D1(n814), .D2(n815), .D3(n812), .D4(n816), .D5(
        n813), .D6(input_log2[40]), .D7(n811), .A(input_log2[45]), .B(
        input_log2[44]), .C(input_log2[43]), .Z(n818) );
  MUX81P U1917 ( .D0(n825), .D1(n822), .D2(n824), .D3(n820), .D4(n284), .D5(
        n821), .D6(n823), .D7(n819), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n826) );
  MUX81P U1918 ( .D0(n834), .D1(n830), .D2(n832), .D3(n828), .D4(n833), .D5(
        n829), .D6(n831), .D7(n827), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n835) );
  MUX81P U1919 ( .D0(n843), .D1(n839), .D2(n841), .D3(n837), .D4(n842), .D5(
        n838), .D6(n840), .D7(n836), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n844) );
  MUX81P U1920 ( .D0(n852), .D1(n848), .D2(n850), .D3(n846), .D4(n851), .D5(
        n847), .D6(n849), .D7(n845), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n853) );
  MUX81P U1921 ( .D0(n868), .D1(n864), .D2(n866), .D3(n862), .D4(n867), .D5(
        n863), .D6(n865), .D7(n861), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n869) );
  MUX81P U1922 ( .D0(n877), .D1(n873), .D2(n875), .D3(n871), .D4(n876), .D5(
        n872), .D6(n874), .D7(n870), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n878) );
  MUX81P U1923 ( .D0(n889), .D1(n885), .D2(n887), .D3(n884), .D4(n888), .D5(
        n234), .D6(n886), .D7(n883), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n890) );
  MUX81P U1924 ( .D0(n897), .D1(n893), .D2(n895), .D3(n891), .D4(n896), .D5(
        n892), .D6(n894), .D7(n224), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n898) );
  MUX81P U1925 ( .D0(n906), .D1(n902), .D2(n904), .D3(n900), .D4(n905), .D5(
        n901), .D6(n903), .D7(n899), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n907) );
  MUX81P U1926 ( .D0(n914), .D1(n911), .D2(n235), .D3(n909), .D4(n913), .D5(
        n910), .D6(n912), .D7(n908), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n915) );
  MUX81P U1927 ( .D0(n923), .D1(n919), .D2(n921), .D3(n917), .D4(n922), .D5(
        n918), .D6(n920), .D7(n916), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n924) );
  MUX81P U1928 ( .D0(n932), .D1(n928), .D2(n930), .D3(n926), .D4(n931), .D5(
        n927), .D6(n929), .D7(n925), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n933) );
  MUX81P U1929 ( .D0(n948), .D1(n944), .D2(n946), .D3(n942), .D4(n947), .D5(
        n943), .D6(n945), .D7(n941), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n949) );
  MUX81P U1930 ( .D0(n957), .D1(n953), .D2(n955), .D3(n951), .D4(n956), .D5(
        n952), .D6(n954), .D7(n950), .A(input_log2[45]), .B(input_log2[44]), 
        .C(input_log2[43]), .Z(n958) );
  AN2P U1931 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n989) );
  AN2P U1932 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n993) );
  AN2P U1933 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n997) );
  AN2P U1934 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1006) );
  AN2P U1935 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1016) );
  AN2P U1936 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1025) );
  AN2P U1937 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1028) );
  AN2P U1938 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1034) );
  AN2P U1939 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1038) );
  AN2P U1940 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1058) );
  AN2P U1941 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1067) );
  AN2P U1942 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1087) );
  AN2P U1943 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1113) );
  AN2P U1944 ( .A(input_log2[42]), .B(input_log2[41]), .Z(n1123) );
  AN2P U1945 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1151) );
  AN2P U1946 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1158) );
  AN2P U1947 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1161) );
  AN2P U1948 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1173) );
  AN2P U1949 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1179) );
  AN2P U1950 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1190) );
  AN2P U1951 ( .A(input_log2[42]), .B(input_log2[40]), .Z(n1195) );
  AN2P U1952 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1204) );
  AN2P U1953 ( .A(input_log2[42]), .B(input_log2[40]), .Z(n1213) );
  AN2P U1954 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1219) );
  AN2P U1955 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1238) );
  AN2P U1956 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1255) );
  AN2P U1957 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1260) );
  AN2P U1958 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1264) );
  AN2P U1959 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1268) );
  AN2P U1960 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1275) );
  AN2P U1961 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1280) );
  AN2P U1962 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1307) );
  AN2P U1963 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1314) );
  AN2P U1964 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1319) );
  AN2P U1965 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1330) );
  AN2P U1966 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1339) );
  AN2P U1967 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1352) );
  AN2P U1968 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1378) );
  AN2P U1969 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1384) );
  AN2P U1970 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1419) );
  AN2P U1971 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1435) );
  AN2P U1972 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1445) );
  AN2P U1973 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1451) );
  AN2P U1974 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1476) );
  AN2P U1975 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1490) );
  AN2P U1976 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1534) );
  AN2P U1977 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1540) );
  AN2P U1978 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1550) );
  AN2P U1979 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1559) );
  AN2P U1980 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1567) );
  AN2P U1981 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1577) );
  AN2P U1982 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1615) );
  AN2P U1983 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1622) );
  AN2P U1984 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1634) );
  AN2P U1985 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1665) );
  AN2P U1986 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1691) );
  AN2P U1987 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1701) );
  AN2P U1988 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1728) );
  AN2P U1989 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1737) );
  AN2P U1990 ( .A(input_log2[40]), .B(input_log2[41]), .Z(n1741) );
  AN2P U1991 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1765) );
  AN2P U1992 ( .A(input_log2[40]), .B(input_log2[42]), .Z(n1784) );
  AN2P U1993 ( .A(input_log2[41]), .B(input_log2[40]), .Z(n1822) );
  AN2P U1994 ( .A(input_log2[41]), .B(input_log2[42]), .Z(n1833) );
  AN2P U1995 ( .A(n630), .B(input_log2[43]), .Z(n1869) );
  AN2P U1996 ( .A(input_log2[43]), .B(n608), .Z(n1876) );
  AN2P U1997 ( .A(input_log2[47]), .B(n295), .Z(n1919) );
  AN2P U1998 ( .A(n348), .B(input_log2[45]), .Z(n1945) );
  AN2P U1999 ( .A(n610), .B(input_log2[45]), .Z(n1955) );
  AN2P U2000 ( .A(input_log2[43]), .B(n593), .Z(n1962) );
  AN2P U2001 ( .A(input_log2[43]), .B(n564), .Z(n2093) );
  AN2P U2002 ( .A(input_log2[43]), .B(input_log2[44]), .Z(n2097) );
  AN2P U2003 ( .A(input_log2[44]), .B(n302), .Z(n2098) );
  AN2P U2004 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n2107) );
  AN2P U2005 ( .A(n767), .B(input_log2[44]), .Z(n2109) );
  AN2P U2006 ( .A(input_log2[44]), .B(n769), .Z(n2111) );
  AN2P U2007 ( .A(input_log2[43]), .B(n768), .Z(n2113) );
  AN2P U2008 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n2119) );
  AN2P U2009 ( .A(n496), .B(input_log2[44]), .Z(n2121) );
  AN2P U2010 ( .A(input_log2[44]), .B(n499), .Z(n2123) );
  AN2P U2011 ( .A(input_log2[43]), .B(n497), .Z(n2125) );
  AN2P U2012 ( .A(n746), .B(input_log2[44]), .Z(n2140) );
  AN2P U2013 ( .A(input_log2[44]), .B(input_log2[45]), .Z(n2183) );
  AN2P U2014 ( .A(n724), .B(input_log2[44]), .Z(n2185) );
  AN2P U2015 ( .A(input_log2[43]), .B(n725), .Z(n2189) );
  AN2P U2016 ( .A(n698), .B(input_log2[44]), .Z(n2196) );
  AN2P U2017 ( .A(n699), .B(input_log2[43]), .Z(n2198) );
  AN2P U2018 ( .A(n225), .B(input_log2[43]), .Z(n2200) );
  IV U2019 ( .A(reset), .Z(n2235) );
  EO U2020 ( .A(n2234), .B(n2216), .Z(N142) );
  NR2 U2021 ( .A(num2_1[66]), .B(n2217), .Z(n2216) );
  EO U2022 ( .A(n2217), .B(num2_1[66]), .Z(N141) );
  ND2 U2023 ( .A(n230), .B(n2218), .Z(n2217) );
  EN U2024 ( .A(num2_1[65]), .B(n2218), .Z(N140) );
  AO4 U2025 ( .A(n2219), .B(n2220), .C(num2_1[64]), .D(n2221), .Z(n2218) );
  AN2 U2026 ( .A(n2220), .B(n2219), .Z(n2221) );
  EN U2027 ( .A(n2219), .B(n2222), .Z(N139) );
  EO U2028 ( .A(n2220), .B(num2_1[64]), .Z(n2222) );
  ND2 U2029 ( .A(num3_1[26]), .B(n2223), .Z(n2220) );
  EO1 U2030 ( .A(n2224), .B(n2225), .C(num2_1[63]), .D(n2226), .Z(n2219) );
  NR2 U2031 ( .A(n2225), .B(n2224), .Z(n2226) );
  EO U2032 ( .A(n2225), .B(n2227), .Z(N138) );
  EN U2033 ( .A(num2_1[63]), .B(n2224), .Z(n2227) );
  EON1 U2034 ( .A(num2_1[62]), .B(n2228), .C(n2229), .D(n2230), .Z(n2224) );
  NR2 U2035 ( .A(n2230), .B(n2229), .Z(n2228) );
  EO U2036 ( .A(n2223), .B(num3_1[26]), .Z(n2225) );
  AN3 U2037 ( .A(num3_1[24]), .B(n229), .C(num3_1[25]), .Z(n2223) );
  EO U2038 ( .A(n2230), .B(n2231), .Z(N137) );
  EN U2039 ( .A(num2_1[62]), .B(n2229), .Z(n2231) );
  EN U2040 ( .A(n2232), .B(num3_1[25]), .Z(n2230) );
  ND2 U2041 ( .A(num3_1[24]), .B(n229), .Z(n2232) );
  AO7 U2042 ( .A(num2_1[61]), .B(n2233), .C(n2229), .Z(N136) );
  ND2 U2043 ( .A(num2_1[61]), .B(n2233), .Z(n2229) );
  EN U2044 ( .A(n229), .B(num3_1[24]), .Z(n2233) );
endmodule


module Poly_sqrt_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;

  wire   [13:1] carry;

  FA1A U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA1A U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA1A U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  FA1A U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA1A U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA1A U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA1A U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA1A U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA1A U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA1A U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA1A U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA1A U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(SUM[13]), .S(SUM[12])
         );
  EO U1 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  AN2P U2 ( .A(A[0]), .B(B[0]), .Z(carry[1]) );
endmodule


module Poly_sqrt_DW01_add_1 ( A, B, CI, SUM, CO );
  input [40:0] A;
  input [40:0] B;
  output [40:0] SUM;
  input CI;
  output CO;
  wire   \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35;
  assign SUM[29] = A[29];
  assign SUM[21] = A[21];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];

  AN2P U2 ( .A(n2), .B(n35), .Z(SUM[30]) );
  IVP U3 ( .A(n26), .Z(n6) );
  IVP U4 ( .A(n18), .Z(n4) );
  IVP U5 ( .A(n33), .Z(n8) );
  IVP U6 ( .A(n20), .Z(n5) );
  IVP U7 ( .A(n12), .Z(n3) );
  IVP U8 ( .A(n28), .Z(n7) );
  IVP U9 ( .A(n35), .Z(n9) );
  OR2 U10 ( .A(B[30]), .B(A[30]), .Z(n2) );
  EO U11 ( .A(n10), .B(n11), .Z(SUM[37]) );
  EO U12 ( .A(B[37]), .B(A[37]), .Z(n11) );
  AO7 U13 ( .A(n12), .B(n13), .C(n14), .Z(n10) );
  EO U14 ( .A(n15), .B(n13), .Z(SUM[36]) );
  AO6 U15 ( .A(n16), .B(n17), .C(n4), .Z(n13) );
  ND2 U16 ( .A(n3), .B(n14), .Z(n15) );
  ND2 U17 ( .A(B[36]), .B(A[36]), .Z(n14) );
  NR2 U18 ( .A(B[36]), .B(A[36]), .Z(n12) );
  EN U19 ( .A(n19), .B(n17), .Z(SUM[35]) );
  AO7 U20 ( .A(n20), .B(n21), .C(n22), .Z(n17) );
  ND2 U21 ( .A(n16), .B(n18), .Z(n19) );
  ND2 U22 ( .A(B[35]), .B(A[35]), .Z(n18) );
  OR2 U23 ( .A(B[35]), .B(A[35]), .Z(n16) );
  EO U24 ( .A(n23), .B(n21), .Z(SUM[34]) );
  AO6 U25 ( .A(n24), .B(n25), .C(n6), .Z(n21) );
  ND2 U26 ( .A(n5), .B(n22), .Z(n23) );
  ND2 U27 ( .A(B[34]), .B(A[34]), .Z(n22) );
  NR2 U28 ( .A(B[34]), .B(A[34]), .Z(n20) );
  EN U29 ( .A(n27), .B(n25), .Z(SUM[33]) );
  AO7 U30 ( .A(n28), .B(n29), .C(n30), .Z(n25) );
  ND2 U31 ( .A(n24), .B(n26), .Z(n27) );
  ND2 U32 ( .A(B[33]), .B(A[33]), .Z(n26) );
  OR2 U33 ( .A(B[33]), .B(A[33]), .Z(n24) );
  EO U34 ( .A(n31), .B(n29), .Z(SUM[32]) );
  AO6 U35 ( .A(n32), .B(n9), .C(n8), .Z(n29) );
  ND2 U36 ( .A(n7), .B(n30), .Z(n31) );
  ND2 U37 ( .A(B[32]), .B(A[32]), .Z(n30) );
  NR2 U38 ( .A(B[32]), .B(A[32]), .Z(n28) );
  EN U39 ( .A(n34), .B(n9), .Z(SUM[31]) );
  ND2 U40 ( .A(n32), .B(n33), .Z(n34) );
  ND2 U41 ( .A(B[31]), .B(A[31]), .Z(n33) );
  OR2 U42 ( .A(B[31]), .B(A[31]), .Z(n32) );
  ND2 U43 ( .A(B[30]), .B(A[30]), .Z(n35) );
endmodule


module Poly_sqrt_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [30:0] A;
  input [11:0] B;
  output [42:0] PRODUCT;
  input TC;
  wire   \ab[30][11] , \ab[30][10] , \ab[30][9] , \ab[30][8] , \ab[30][7] ,
         \ab[30][6] , \ab[30][5] , \ab[30][4] , \ab[30][3] , \ab[30][2] ,
         \ab[30][1] , \ab[30][0] , \ab[29][11] , \ab[29][10] , \ab[29][9] ,
         \ab[29][8] , \ab[29][7] , \ab[29][6] , \ab[29][5] , \ab[29][4] ,
         \ab[29][3] , \ab[29][2] , \ab[29][1] , \ab[29][0] , \ab[28][11] ,
         \ab[28][10] , \ab[28][9] , \ab[28][8] , \ab[28][7] , \ab[28][6] ,
         \ab[28][5] , \ab[28][4] , \ab[28][3] , \ab[28][2] , \ab[28][1] ,
         \ab[28][0] , \ab[27][11] , \ab[27][10] , \ab[27][9] , \ab[27][8] ,
         \ab[27][7] , \ab[27][6] , \ab[27][5] , \ab[27][4] , \ab[27][3] ,
         \ab[27][2] , \ab[27][1] , \ab[27][0] , \ab[26][11] , \ab[26][10] ,
         \ab[26][9] , \ab[26][8] , \ab[26][7] , \ab[26][6] , \ab[26][5] ,
         \ab[26][4] , \ab[26][3] , \ab[26][2] , \ab[26][1] , \ab[26][0] ,
         \ab[25][11] , \ab[25][10] , \ab[25][9] , \ab[25][8] , \ab[25][7] ,
         \ab[25][6] , \ab[25][5] , \ab[25][4] , \ab[25][3] , \ab[25][2] ,
         \ab[25][1] , \ab[25][0] , \ab[24][11] , \ab[24][10] , \ab[24][9] ,
         \ab[24][8] , \ab[24][7] , \ab[24][6] , \ab[24][5] , \ab[24][4] ,
         \ab[24][3] , \ab[24][2] , \ab[24][1] , \ab[24][0] , \ab[23][11] ,
         \ab[23][10] , \ab[23][9] , \ab[23][8] , \ab[23][7] , \ab[23][6] ,
         \ab[23][5] , \ab[23][4] , \ab[23][3] , \ab[23][2] , \ab[23][1] ,
         \ab[23][0] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][11] , \ab[21][10] ,
         \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] , \ab[21][5] ,
         \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] ,
         \ab[20][11] , \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] ,
         \ab[20][6] , \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] ,
         \ab[20][1] , \ab[20][0] , \ab[19][11] , \ab[19][10] , \ab[19][9] ,
         \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] ,
         \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][11] ,
         \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] , \ab[18][6] ,
         \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] , \ab[18][1] ,
         \ab[18][0] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][11] , \ab[16][10] ,
         \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] , \ab[16][5] ,
         \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] , \ab[16][0] ,
         \ab[15][11] , \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] ,
         \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] ,
         \ab[15][1] , \ab[15][0] , \ab[14][11] , \ab[14][10] , \ab[14][9] ,
         \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] ,
         \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][11] ,
         \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] , \ab[13][6] ,
         \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] , \ab[13][1] ,
         \ab[13][0] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] ,
         \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] ,
         \ab[10][1] , \ab[10][0] , \ab[9][11] , \ab[9][10] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][11] ,
         \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] ,
         \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] ,
         \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] ,
         \ab[5][1] , \ab[5][0] , \ab[4][11] , \ab[4][10] , \ab[4][9] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[30][10] ,
         \CARRYB[30][9] , \CARRYB[30][8] , \CARRYB[30][7] , \CARRYB[30][6] ,
         \CARRYB[30][5] , \CARRYB[30][4] , \CARRYB[30][3] , \CARRYB[30][2] ,
         \CARRYB[30][1] , \CARRYB[30][0] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][10] , \CARRYB[28][9] , \CARRYB[28][8] ,
         \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] , \CARRYB[28][4] ,
         \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] ,
         \CARRYB[27][10] , \CARRYB[27][9] , \CARRYB[27][8] , \CARRYB[27][7] ,
         \CARRYB[27][6] , \CARRYB[27][5] , \CARRYB[27][4] , \CARRYB[27][3] ,
         \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] , \CARRYB[26][10] ,
         \CARRYB[26][9] , \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] ,
         \CARRYB[26][5] , \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] ,
         \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][10] , \CARRYB[25][9] ,
         \CARRYB[25][8] , \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][10] , \CARRYB[24][9] , \CARRYB[24][8] ,
         \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] ,
         \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] , \CARRYB[23][7] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][10] ,
         \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] ,
         \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] ,
         \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] ,
         \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][10] ,
         \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] ,
         \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] ,
         \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] ,
         \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] ,
         \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][10] ,
         \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] ,
         \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] ,
         \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][10] ,
         \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][10] ,
         \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][10] ,
         \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[30][10] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[30][0] ,
         \SUMB[29][10] , \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] ,
         \SUMB[29][6] , \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] ,
         \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][10] , \SUMB[28][9] ,
         \SUMB[28][8] , \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] ,
         \SUMB[28][4] , \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] ,
         \SUMB[27][10] , \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] ,
         \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][10] , \SUMB[26][9] ,
         \SUMB[26][8] , \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] ,
         \SUMB[26][4] , \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] ,
         \SUMB[25][10] , \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][10] , \SUMB[24][9] ,
         \SUMB[24][8] , \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] ,
         \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][10] , \SUMB[22][9] ,
         \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] ,
         \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][10] , \SUMB[20][9] ,
         \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] ,
         \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][10] , \SUMB[18][9] ,
         \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] ,
         \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] ,
         \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] ,
         \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] ,
         \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][10] , \SUMB[16][9] ,
         \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \PROD1[11] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] ,
         \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[27] ,
         \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] ,
         \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] ,
         \A1[12] , \A1[11] , \A1[10] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[40] , \A2[39] ,
         \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] ,
         \A2[31] , \A2[30] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  Poly_sqrt_DW01_add_1 FS_1 ( .A({1'b0, \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \SUMB[30][0] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , 
        \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \PROD1[11] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , 
        \A1[2] , \A1[1] , \A1[0] }), .B({\A2[40] , \A2[39] , \A2[38] , 
        \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , 
        \A2[30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, PRODUCT[39:23], SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S5_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\ab[29][11] ), .CO(
        \CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA1A S4_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), .CO(
        \CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA1A S4_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), .CO(
        \CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA1A S3_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\ab[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA1A S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA1A S3_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\ab[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA1A S4_3 ( .A(\ab[30][3] ), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), .CO(
        \CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA1A S4_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), .CO(
        \CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA1A S4_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), .CO(
        \CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA1A S4_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), .CO(
        \CARRYB[30][0] ), .S(\SUMB[30][0] ) );
  FA1A S4_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), .CO(
        \CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA1A S4_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), .CO(
        \CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA1A S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA1A S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA1A S2_29_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA1A S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FA1A S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA1A S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA1A S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA1A S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA1A S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA1A S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA1A S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA1A S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA1A S3_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\ab[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA1A S4_4 ( .A(\ab[30][4] ), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), .CO(
        \CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA1A S4_5 ( .A(\ab[30][5] ), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), .CO(
        \CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA1A S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA1A S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA1A S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA1A S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA1A S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA1A S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA1A S2_29_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA1A S2_29_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA1A S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA1A S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA1A S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA1A S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA1A S3_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\ab[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA1A S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA1A S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA1A S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA1A S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA1A S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA1A S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA1A S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA1A S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA1A S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA1A S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA1A S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA1A S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA1A S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA1A S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA1A S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA1A S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA1A S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA1A S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA1A S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA1A S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA1A S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA1A S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA1A S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA1A S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA1A S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA1A S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA1A S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA1A S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA1A S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA1A S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA1A S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA1A S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA1A S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA1A S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA1A S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA1A S3_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\ab[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA1A S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA1A S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA1A S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA1A S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA1A S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA1A S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA1A S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA1A S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA1A S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA1A S3_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\ab[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA1A S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA1A S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA1A S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA1A S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA1A S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA1A S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA1A S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA1A S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA1A S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA1A S3_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\ab[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA1A S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA1A S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA1A S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA1A S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA1A S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA1A S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA1A S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA1A S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA1A S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA1A S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA1A S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA1A S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA1A S3_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\ab[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA1A S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA1A S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA1A S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA1A S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA1A S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA1A S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA1A S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA1A S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA1A S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA1A S3_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\ab[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA1A S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA1A S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA1A S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA1A S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA1A S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA1A S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA1A S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA1A S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA1A S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA1A S3_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\ab[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA1A S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA1A S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA1A S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA1A S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA1A S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA1A S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA1A S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA1A S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA1A S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA1A S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA1A S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA1A S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA1A S3_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\ab[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA1A S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA1A S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA1A S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA1A S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA1A S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA1A S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA1A S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA1A S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA1A S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA1A S3_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\ab[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA1A S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA1A S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA1A S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA1A S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA1A S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA1A S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA1A S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA1A S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA1A S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA1A S3_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\ab[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA1A S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA1A S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA1A S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA1A S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA1A S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA1A S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA1A S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA1A S3_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\ab[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA1A S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA1A S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA1A S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA1A S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA1A S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA1A S3_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\ab[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S3_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\ab[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\PROD1[11] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S3_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\ab[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S3_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\ab[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S3_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\ab[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S3_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\ab[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S3_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\ab[8][11] ), .CO(
        \CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S3_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\ab[7][11] ), .CO(
        \CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S3_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\ab[6][11] ), .CO(
        \CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S3_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\ab[5][11] ), .CO(
        \CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S3_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\ab[4][11] ), .CO(
        \CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S3_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\ab[3][11] ), .CO(
        \CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S3_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\ab[2][11] ), .CO(
        \CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S3_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\ab[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  EO U2 ( .A(\CARRYB[30][8] ), .B(\SUMB[30][9] ), .Z(\A1[37] ) );
  EO U3 ( .A(\CARRYB[30][5] ), .B(\SUMB[30][6] ), .Z(\A1[34] ) );
  EO U4 ( .A(\CARRYB[30][7] ), .B(\SUMB[30][8] ), .Z(\A1[36] ) );
  EO U5 ( .A(\CARRYB[30][1] ), .B(\SUMB[30][2] ), .Z(\A1[30] ) );
  EO U6 ( .A(\CARRYB[30][3] ), .B(\SUMB[30][4] ), .Z(\A1[32] ) );
  EO U7 ( .A(\CARRYB[30][6] ), .B(\SUMB[30][7] ), .Z(\A1[35] ) );
  EO U8 ( .A(\CARRYB[30][2] ), .B(\SUMB[30][3] ), .Z(\A1[31] ) );
  EO U9 ( .A(\CARRYB[30][4] ), .B(\SUMB[30][5] ), .Z(\A1[33] ) );
  EO U10 ( .A(\CARRYB[30][9] ), .B(\SUMB[30][10] ), .Z(\A1[38] ) );
  EO U11 ( .A(\CARRYB[30][10] ), .B(\ab[30][11] ), .Z(\A1[39] ) );
  IVP U12 ( .A(B[10]), .Z(n10) );
  IVP U13 ( .A(B[9]), .Z(n9) );
  IVP U14 ( .A(B[0]), .Z(n12) );
  EO U15 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U16 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U17 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U18 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U19 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U20 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U21 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  EO U22 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U23 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  IVP U24 ( .A(B[8]), .Z(n8) );
  IVP U25 ( .A(B[7]), .Z(n15) );
  IVP U26 ( .A(B[6]), .Z(n14) );
  IVP U27 ( .A(B[5]), .Z(n13) );
  IVP U28 ( .A(B[4]), .Z(n4) );
  IVP U29 ( .A(B[11]), .Z(n11) );
  IVP U30 ( .A(B[3]), .Z(n5) );
  IVP U31 ( .A(B[2]), .Z(n6) );
  IVP U32 ( .A(B[1]), .Z(n7) );
  IVP U33 ( .A(A[3]), .Z(n42) );
  IVP U34 ( .A(A[2]), .Z(n43) );
  IVP U35 ( .A(A[4]), .Z(n41) );
  IVP U36 ( .A(A[6]), .Z(n39) );
  IVP U37 ( .A(A[5]), .Z(n40) );
  IVP U38 ( .A(A[7]), .Z(n38) );
  IVP U39 ( .A(A[9]), .Z(n36) );
  IVP U40 ( .A(A[8]), .Z(n37) );
  IVP U41 ( .A(A[10]), .Z(n35) );
  IVP U42 ( .A(A[12]), .Z(n33) );
  IVP U43 ( .A(A[11]), .Z(n34) );
  IVP U44 ( .A(A[13]), .Z(n32) );
  IVP U45 ( .A(A[15]), .Z(n30) );
  IVP U46 ( .A(A[14]), .Z(n31) );
  IVP U47 ( .A(A[16]), .Z(n29) );
  IVP U48 ( .A(A[18]), .Z(n27) );
  IVP U49 ( .A(A[17]), .Z(n28) );
  IVP U50 ( .A(A[19]), .Z(n26) );
  IVP U51 ( .A(A[21]), .Z(n24) );
  IVP U52 ( .A(A[20]), .Z(n25) );
  IVP U53 ( .A(A[22]), .Z(n23) );
  IVP U54 ( .A(A[24]), .Z(n21) );
  IVP U55 ( .A(A[25]), .Z(n20) );
  IVP U56 ( .A(A[23]), .Z(n22) );
  IVP U57 ( .A(A[26]), .Z(n19) );
  IVP U58 ( .A(A[27]), .Z(n18) );
  IVP U59 ( .A(A[28]), .Z(n17) );
  IVP U60 ( .A(A[29]), .Z(n16) );
  IVP U61 ( .A(A[30]), .Z(n3) );
  IVP U62 ( .A(A[1]), .Z(n44) );
  EO U63 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  EO U64 ( .A(\CARRYB[30][0] ), .B(\SUMB[30][1] ), .Z(\A1[29] ) );
  IVP U65 ( .A(A[0]), .Z(n45) );
  AN2P U66 ( .A(\CARRYB[30][0] ), .B(\SUMB[30][1] ), .Z(\A2[30] ) );
  AN2P U67 ( .A(\CARRYB[30][1] ), .B(\SUMB[30][2] ), .Z(\A2[31] ) );
  AN2P U68 ( .A(\CARRYB[30][2] ), .B(\SUMB[30][3] ), .Z(\A2[32] ) );
  AN2P U69 ( .A(\CARRYB[30][3] ), .B(\SUMB[30][4] ), .Z(\A2[33] ) );
  AN2P U70 ( .A(\CARRYB[30][4] ), .B(\SUMB[30][5] ), .Z(\A2[34] ) );
  AN2P U71 ( .A(\CARRYB[30][5] ), .B(\SUMB[30][6] ), .Z(\A2[35] ) );
  AN2P U72 ( .A(\CARRYB[30][6] ), .B(\SUMB[30][7] ), .Z(\A2[36] ) );
  AN2P U73 ( .A(\CARRYB[30][7] ), .B(\SUMB[30][8] ), .Z(\A2[37] ) );
  AN2P U74 ( .A(\CARRYB[30][8] ), .B(\SUMB[30][9] ), .Z(\A2[38] ) );
  AN2P U75 ( .A(\CARRYB[30][9] ), .B(\SUMB[30][10] ), .Z(\A2[39] ) );
  AN2P U76 ( .A(\CARRYB[30][10] ), .B(\ab[30][11] ), .Z(\A2[40] ) );
  AN2P U77 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U78 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U79 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U80 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U81 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U82 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U83 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U84 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U85 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U86 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  NR2 U88 ( .A(n36), .B(n9), .Z(\ab[9][9] ) );
  NR2 U89 ( .A(n36), .B(n8), .Z(\ab[9][8] ) );
  NR2 U90 ( .A(n36), .B(n15), .Z(\ab[9][7] ) );
  NR2 U91 ( .A(n36), .B(n14), .Z(\ab[9][6] ) );
  NR2 U92 ( .A(n36), .B(n13), .Z(\ab[9][5] ) );
  NR2 U93 ( .A(n36), .B(n4), .Z(\ab[9][4] ) );
  NR2 U94 ( .A(n36), .B(n5), .Z(\ab[9][3] ) );
  NR2 U95 ( .A(n36), .B(n6), .Z(\ab[9][2] ) );
  NR2 U96 ( .A(n36), .B(n7), .Z(\ab[9][1] ) );
  NR2 U97 ( .A(n36), .B(n11), .Z(\ab[9][11] ) );
  NR2 U98 ( .A(n36), .B(n10), .Z(\ab[9][10] ) );
  NR2 U99 ( .A(n36), .B(n12), .Z(\ab[9][0] ) );
  NR2 U100 ( .A(n9), .B(n37), .Z(\ab[8][9] ) );
  NR2 U101 ( .A(n8), .B(n37), .Z(\ab[8][8] ) );
  NR2 U102 ( .A(n15), .B(n37), .Z(\ab[8][7] ) );
  NR2 U103 ( .A(n14), .B(n37), .Z(\ab[8][6] ) );
  NR2 U104 ( .A(n13), .B(n37), .Z(\ab[8][5] ) );
  NR2 U105 ( .A(n4), .B(n37), .Z(\ab[8][4] ) );
  NR2 U106 ( .A(n5), .B(n37), .Z(\ab[8][3] ) );
  NR2 U107 ( .A(n6), .B(n37), .Z(\ab[8][2] ) );
  NR2 U108 ( .A(n7), .B(n37), .Z(\ab[8][1] ) );
  NR2 U109 ( .A(n11), .B(n37), .Z(\ab[8][11] ) );
  NR2 U110 ( .A(n10), .B(n37), .Z(\ab[8][10] ) );
  NR2 U111 ( .A(n12), .B(n37), .Z(\ab[8][0] ) );
  NR2 U112 ( .A(n9), .B(n38), .Z(\ab[7][9] ) );
  NR2 U113 ( .A(n8), .B(n38), .Z(\ab[7][8] ) );
  NR2 U114 ( .A(n15), .B(n38), .Z(\ab[7][7] ) );
  NR2 U115 ( .A(n14), .B(n38), .Z(\ab[7][6] ) );
  NR2 U116 ( .A(n13), .B(n38), .Z(\ab[7][5] ) );
  NR2 U117 ( .A(n4), .B(n38), .Z(\ab[7][4] ) );
  NR2 U118 ( .A(n5), .B(n38), .Z(\ab[7][3] ) );
  NR2 U119 ( .A(n6), .B(n38), .Z(\ab[7][2] ) );
  NR2 U120 ( .A(n7), .B(n38), .Z(\ab[7][1] ) );
  NR2 U121 ( .A(n11), .B(n38), .Z(\ab[7][11] ) );
  NR2 U122 ( .A(n10), .B(n38), .Z(\ab[7][10] ) );
  NR2 U123 ( .A(n12), .B(n38), .Z(\ab[7][0] ) );
  NR2 U124 ( .A(n9), .B(n39), .Z(\ab[6][9] ) );
  NR2 U125 ( .A(n8), .B(n39), .Z(\ab[6][8] ) );
  NR2 U126 ( .A(n15), .B(n39), .Z(\ab[6][7] ) );
  NR2 U127 ( .A(n14), .B(n39), .Z(\ab[6][6] ) );
  NR2 U128 ( .A(n13), .B(n39), .Z(\ab[6][5] ) );
  NR2 U129 ( .A(n4), .B(n39), .Z(\ab[6][4] ) );
  NR2 U130 ( .A(n5), .B(n39), .Z(\ab[6][3] ) );
  NR2 U131 ( .A(n6), .B(n39), .Z(\ab[6][2] ) );
  NR2 U132 ( .A(n7), .B(n39), .Z(\ab[6][1] ) );
  NR2 U133 ( .A(n11), .B(n39), .Z(\ab[6][11] ) );
  NR2 U134 ( .A(n10), .B(n39), .Z(\ab[6][10] ) );
  NR2 U135 ( .A(n12), .B(n39), .Z(\ab[6][0] ) );
  NR2 U136 ( .A(n9), .B(n40), .Z(\ab[5][9] ) );
  NR2 U137 ( .A(n8), .B(n40), .Z(\ab[5][8] ) );
  NR2 U138 ( .A(n15), .B(n40), .Z(\ab[5][7] ) );
  NR2 U139 ( .A(n14), .B(n40), .Z(\ab[5][6] ) );
  NR2 U140 ( .A(n13), .B(n40), .Z(\ab[5][5] ) );
  NR2 U141 ( .A(n4), .B(n40), .Z(\ab[5][4] ) );
  NR2 U142 ( .A(n5), .B(n40), .Z(\ab[5][3] ) );
  NR2 U143 ( .A(n6), .B(n40), .Z(\ab[5][2] ) );
  NR2 U144 ( .A(n7), .B(n40), .Z(\ab[5][1] ) );
  NR2 U145 ( .A(n11), .B(n40), .Z(\ab[5][11] ) );
  NR2 U146 ( .A(n10), .B(n40), .Z(\ab[5][10] ) );
  NR2 U147 ( .A(n12), .B(n40), .Z(\ab[5][0] ) );
  NR2 U148 ( .A(n9), .B(n41), .Z(\ab[4][9] ) );
  NR2 U149 ( .A(n8), .B(n41), .Z(\ab[4][8] ) );
  NR2 U150 ( .A(n15), .B(n41), .Z(\ab[4][7] ) );
  NR2 U151 ( .A(n14), .B(n41), .Z(\ab[4][6] ) );
  NR2 U152 ( .A(n13), .B(n41), .Z(\ab[4][5] ) );
  NR2 U153 ( .A(n4), .B(n41), .Z(\ab[4][4] ) );
  NR2 U154 ( .A(n5), .B(n41), .Z(\ab[4][3] ) );
  NR2 U155 ( .A(n6), .B(n41), .Z(\ab[4][2] ) );
  NR2 U156 ( .A(n7), .B(n41), .Z(\ab[4][1] ) );
  NR2 U157 ( .A(n11), .B(n41), .Z(\ab[4][11] ) );
  NR2 U158 ( .A(n10), .B(n41), .Z(\ab[4][10] ) );
  NR2 U159 ( .A(n12), .B(n41), .Z(\ab[4][0] ) );
  NR2 U160 ( .A(n9), .B(n42), .Z(\ab[3][9] ) );
  NR2 U161 ( .A(n8), .B(n42), .Z(\ab[3][8] ) );
  NR2 U162 ( .A(n15), .B(n42), .Z(\ab[3][7] ) );
  NR2 U163 ( .A(n14), .B(n42), .Z(\ab[3][6] ) );
  NR2 U164 ( .A(n13), .B(n42), .Z(\ab[3][5] ) );
  NR2 U165 ( .A(n4), .B(n42), .Z(\ab[3][4] ) );
  NR2 U166 ( .A(n5), .B(n42), .Z(\ab[3][3] ) );
  NR2 U167 ( .A(n6), .B(n42), .Z(\ab[3][2] ) );
  NR2 U168 ( .A(n7), .B(n42), .Z(\ab[3][1] ) );
  NR2 U169 ( .A(n11), .B(n42), .Z(\ab[3][11] ) );
  NR2 U170 ( .A(n10), .B(n42), .Z(\ab[3][10] ) );
  NR2 U171 ( .A(n12), .B(n42), .Z(\ab[3][0] ) );
  NR2 U172 ( .A(n9), .B(n3), .Z(\ab[30][9] ) );
  NR2 U173 ( .A(n8), .B(n3), .Z(\ab[30][8] ) );
  NR2 U174 ( .A(n15), .B(n3), .Z(\ab[30][7] ) );
  NR2 U175 ( .A(n14), .B(n3), .Z(\ab[30][6] ) );
  NR2 U176 ( .A(n13), .B(n3), .Z(\ab[30][5] ) );
  NR2 U177 ( .A(n4), .B(n3), .Z(\ab[30][4] ) );
  NR2 U178 ( .A(n5), .B(n3), .Z(\ab[30][3] ) );
  NR2 U179 ( .A(n6), .B(n3), .Z(\ab[30][2] ) );
  NR2 U180 ( .A(n7), .B(n3), .Z(\ab[30][1] ) );
  NR2 U181 ( .A(n11), .B(n3), .Z(\ab[30][11] ) );
  NR2 U182 ( .A(n10), .B(n3), .Z(\ab[30][10] ) );
  NR2 U183 ( .A(n12), .B(n3), .Z(\ab[30][0] ) );
  NR2 U184 ( .A(n9), .B(n43), .Z(\ab[2][9] ) );
  NR2 U185 ( .A(n8), .B(n43), .Z(\ab[2][8] ) );
  NR2 U186 ( .A(n15), .B(n43), .Z(\ab[2][7] ) );
  NR2 U187 ( .A(n14), .B(n43), .Z(\ab[2][6] ) );
  NR2 U188 ( .A(n13), .B(n43), .Z(\ab[2][5] ) );
  NR2 U189 ( .A(n4), .B(n43), .Z(\ab[2][4] ) );
  NR2 U190 ( .A(n5), .B(n43), .Z(\ab[2][3] ) );
  NR2 U191 ( .A(n6), .B(n43), .Z(\ab[2][2] ) );
  NR2 U192 ( .A(n7), .B(n43), .Z(\ab[2][1] ) );
  NR2 U193 ( .A(n11), .B(n43), .Z(\ab[2][11] ) );
  NR2 U194 ( .A(n10), .B(n43), .Z(\ab[2][10] ) );
  NR2 U195 ( .A(n12), .B(n43), .Z(\ab[2][0] ) );
  NR2 U196 ( .A(n9), .B(n16), .Z(\ab[29][9] ) );
  NR2 U197 ( .A(n8), .B(n16), .Z(\ab[29][8] ) );
  NR2 U198 ( .A(n15), .B(n16), .Z(\ab[29][7] ) );
  NR2 U199 ( .A(n14), .B(n16), .Z(\ab[29][6] ) );
  NR2 U200 ( .A(n13), .B(n16), .Z(\ab[29][5] ) );
  NR2 U201 ( .A(n4), .B(n16), .Z(\ab[29][4] ) );
  NR2 U202 ( .A(n5), .B(n16), .Z(\ab[29][3] ) );
  NR2 U203 ( .A(n6), .B(n16), .Z(\ab[29][2] ) );
  NR2 U204 ( .A(n7), .B(n16), .Z(\ab[29][1] ) );
  NR2 U205 ( .A(n11), .B(n16), .Z(\ab[29][11] ) );
  NR2 U206 ( .A(n10), .B(n16), .Z(\ab[29][10] ) );
  NR2 U207 ( .A(n12), .B(n16), .Z(\ab[29][0] ) );
  NR2 U208 ( .A(n9), .B(n17), .Z(\ab[28][9] ) );
  NR2 U209 ( .A(n8), .B(n17), .Z(\ab[28][8] ) );
  NR2 U210 ( .A(n15), .B(n17), .Z(\ab[28][7] ) );
  NR2 U211 ( .A(n14), .B(n17), .Z(\ab[28][6] ) );
  NR2 U212 ( .A(n13), .B(n17), .Z(\ab[28][5] ) );
  NR2 U213 ( .A(n4), .B(n17), .Z(\ab[28][4] ) );
  NR2 U214 ( .A(n5), .B(n17), .Z(\ab[28][3] ) );
  NR2 U215 ( .A(n6), .B(n17), .Z(\ab[28][2] ) );
  NR2 U216 ( .A(n7), .B(n17), .Z(\ab[28][1] ) );
  NR2 U217 ( .A(n11), .B(n17), .Z(\ab[28][11] ) );
  NR2 U218 ( .A(n10), .B(n17), .Z(\ab[28][10] ) );
  NR2 U219 ( .A(n12), .B(n17), .Z(\ab[28][0] ) );
  NR2 U220 ( .A(n9), .B(n18), .Z(\ab[27][9] ) );
  NR2 U221 ( .A(n8), .B(n18), .Z(\ab[27][8] ) );
  NR2 U222 ( .A(n15), .B(n18), .Z(\ab[27][7] ) );
  NR2 U223 ( .A(n14), .B(n18), .Z(\ab[27][6] ) );
  NR2 U224 ( .A(n13), .B(n18), .Z(\ab[27][5] ) );
  NR2 U225 ( .A(n4), .B(n18), .Z(\ab[27][4] ) );
  NR2 U226 ( .A(n5), .B(n18), .Z(\ab[27][3] ) );
  NR2 U227 ( .A(n6), .B(n18), .Z(\ab[27][2] ) );
  NR2 U228 ( .A(n7), .B(n18), .Z(\ab[27][1] ) );
  NR2 U229 ( .A(n11), .B(n18), .Z(\ab[27][11] ) );
  NR2 U230 ( .A(n10), .B(n18), .Z(\ab[27][10] ) );
  NR2 U231 ( .A(n12), .B(n18), .Z(\ab[27][0] ) );
  NR2 U232 ( .A(n9), .B(n19), .Z(\ab[26][9] ) );
  NR2 U233 ( .A(n8), .B(n19), .Z(\ab[26][8] ) );
  NR2 U234 ( .A(n15), .B(n19), .Z(\ab[26][7] ) );
  NR2 U235 ( .A(n14), .B(n19), .Z(\ab[26][6] ) );
  NR2 U236 ( .A(n13), .B(n19), .Z(\ab[26][5] ) );
  NR2 U237 ( .A(n4), .B(n19), .Z(\ab[26][4] ) );
  NR2 U238 ( .A(n5), .B(n19), .Z(\ab[26][3] ) );
  NR2 U239 ( .A(n6), .B(n19), .Z(\ab[26][2] ) );
  NR2 U240 ( .A(n7), .B(n19), .Z(\ab[26][1] ) );
  NR2 U241 ( .A(n11), .B(n19), .Z(\ab[26][11] ) );
  NR2 U242 ( .A(n10), .B(n19), .Z(\ab[26][10] ) );
  NR2 U243 ( .A(n12), .B(n19), .Z(\ab[26][0] ) );
  NR2 U244 ( .A(n9), .B(n20), .Z(\ab[25][9] ) );
  NR2 U245 ( .A(n8), .B(n20), .Z(\ab[25][8] ) );
  NR2 U246 ( .A(n15), .B(n20), .Z(\ab[25][7] ) );
  NR2 U247 ( .A(n14), .B(n20), .Z(\ab[25][6] ) );
  NR2 U248 ( .A(n13), .B(n20), .Z(\ab[25][5] ) );
  NR2 U249 ( .A(n4), .B(n20), .Z(\ab[25][4] ) );
  NR2 U250 ( .A(n5), .B(n20), .Z(\ab[25][3] ) );
  NR2 U251 ( .A(n6), .B(n20), .Z(\ab[25][2] ) );
  NR2 U252 ( .A(n7), .B(n20), .Z(\ab[25][1] ) );
  NR2 U253 ( .A(n11), .B(n20), .Z(\ab[25][11] ) );
  NR2 U254 ( .A(n10), .B(n20), .Z(\ab[25][10] ) );
  NR2 U255 ( .A(n12), .B(n20), .Z(\ab[25][0] ) );
  NR2 U256 ( .A(n9), .B(n21), .Z(\ab[24][9] ) );
  NR2 U257 ( .A(n8), .B(n21), .Z(\ab[24][8] ) );
  NR2 U258 ( .A(n15), .B(n21), .Z(\ab[24][7] ) );
  NR2 U259 ( .A(n14), .B(n21), .Z(\ab[24][6] ) );
  NR2 U260 ( .A(n13), .B(n21), .Z(\ab[24][5] ) );
  NR2 U261 ( .A(n4), .B(n21), .Z(\ab[24][4] ) );
  NR2 U262 ( .A(n5), .B(n21), .Z(\ab[24][3] ) );
  NR2 U263 ( .A(n6), .B(n21), .Z(\ab[24][2] ) );
  NR2 U264 ( .A(n7), .B(n21), .Z(\ab[24][1] ) );
  NR2 U265 ( .A(n11), .B(n21), .Z(\ab[24][11] ) );
  NR2 U266 ( .A(n10), .B(n21), .Z(\ab[24][10] ) );
  NR2 U267 ( .A(n12), .B(n21), .Z(\ab[24][0] ) );
  NR2 U268 ( .A(n9), .B(n22), .Z(\ab[23][9] ) );
  NR2 U269 ( .A(n8), .B(n22), .Z(\ab[23][8] ) );
  NR2 U270 ( .A(n15), .B(n22), .Z(\ab[23][7] ) );
  NR2 U271 ( .A(n14), .B(n22), .Z(\ab[23][6] ) );
  NR2 U272 ( .A(n13), .B(n22), .Z(\ab[23][5] ) );
  NR2 U273 ( .A(n4), .B(n22), .Z(\ab[23][4] ) );
  NR2 U274 ( .A(n5), .B(n22), .Z(\ab[23][3] ) );
  NR2 U275 ( .A(n6), .B(n22), .Z(\ab[23][2] ) );
  NR2 U276 ( .A(n7), .B(n22), .Z(\ab[23][1] ) );
  NR2 U277 ( .A(n11), .B(n22), .Z(\ab[23][11] ) );
  NR2 U278 ( .A(n10), .B(n22), .Z(\ab[23][10] ) );
  NR2 U279 ( .A(n12), .B(n22), .Z(\ab[23][0] ) );
  NR2 U280 ( .A(n9), .B(n23), .Z(\ab[22][9] ) );
  NR2 U281 ( .A(n8), .B(n23), .Z(\ab[22][8] ) );
  NR2 U282 ( .A(n15), .B(n23), .Z(\ab[22][7] ) );
  NR2 U283 ( .A(n14), .B(n23), .Z(\ab[22][6] ) );
  NR2 U284 ( .A(n13), .B(n23), .Z(\ab[22][5] ) );
  NR2 U285 ( .A(n4), .B(n23), .Z(\ab[22][4] ) );
  NR2 U286 ( .A(n5), .B(n23), .Z(\ab[22][3] ) );
  NR2 U287 ( .A(n6), .B(n23), .Z(\ab[22][2] ) );
  NR2 U288 ( .A(n7), .B(n23), .Z(\ab[22][1] ) );
  NR2 U289 ( .A(n11), .B(n23), .Z(\ab[22][11] ) );
  NR2 U290 ( .A(n10), .B(n23), .Z(\ab[22][10] ) );
  NR2 U291 ( .A(n12), .B(n23), .Z(\ab[22][0] ) );
  NR2 U292 ( .A(n9), .B(n24), .Z(\ab[21][9] ) );
  NR2 U293 ( .A(n8), .B(n24), .Z(\ab[21][8] ) );
  NR2 U294 ( .A(n15), .B(n24), .Z(\ab[21][7] ) );
  NR2 U295 ( .A(n14), .B(n24), .Z(\ab[21][6] ) );
  NR2 U296 ( .A(n13), .B(n24), .Z(\ab[21][5] ) );
  NR2 U297 ( .A(n4), .B(n24), .Z(\ab[21][4] ) );
  NR2 U298 ( .A(n5), .B(n24), .Z(\ab[21][3] ) );
  NR2 U299 ( .A(n6), .B(n24), .Z(\ab[21][2] ) );
  NR2 U300 ( .A(n7), .B(n24), .Z(\ab[21][1] ) );
  NR2 U301 ( .A(n11), .B(n24), .Z(\ab[21][11] ) );
  NR2 U302 ( .A(n10), .B(n24), .Z(\ab[21][10] ) );
  NR2 U303 ( .A(n12), .B(n24), .Z(\ab[21][0] ) );
  NR2 U304 ( .A(n9), .B(n25), .Z(\ab[20][9] ) );
  NR2 U305 ( .A(n8), .B(n25), .Z(\ab[20][8] ) );
  NR2 U306 ( .A(n15), .B(n25), .Z(\ab[20][7] ) );
  NR2 U307 ( .A(n14), .B(n25), .Z(\ab[20][6] ) );
  NR2 U308 ( .A(n13), .B(n25), .Z(\ab[20][5] ) );
  NR2 U309 ( .A(n4), .B(n25), .Z(\ab[20][4] ) );
  NR2 U310 ( .A(n5), .B(n25), .Z(\ab[20][3] ) );
  NR2 U311 ( .A(n6), .B(n25), .Z(\ab[20][2] ) );
  NR2 U312 ( .A(n7), .B(n25), .Z(\ab[20][1] ) );
  NR2 U313 ( .A(n11), .B(n25), .Z(\ab[20][11] ) );
  NR2 U314 ( .A(n10), .B(n25), .Z(\ab[20][10] ) );
  NR2 U315 ( .A(n12), .B(n25), .Z(\ab[20][0] ) );
  NR2 U316 ( .A(n9), .B(n44), .Z(\ab[1][9] ) );
  NR2 U317 ( .A(n8), .B(n44), .Z(\ab[1][8] ) );
  NR2 U318 ( .A(n15), .B(n44), .Z(\ab[1][7] ) );
  NR2 U319 ( .A(n14), .B(n44), .Z(\ab[1][6] ) );
  NR2 U320 ( .A(n13), .B(n44), .Z(\ab[1][5] ) );
  NR2 U321 ( .A(n4), .B(n44), .Z(\ab[1][4] ) );
  NR2 U322 ( .A(n5), .B(n44), .Z(\ab[1][3] ) );
  NR2 U323 ( .A(n6), .B(n44), .Z(\ab[1][2] ) );
  NR2 U324 ( .A(n11), .B(n44), .Z(\ab[1][11] ) );
  NR2 U325 ( .A(n10), .B(n44), .Z(\ab[1][10] ) );
  NR2 U326 ( .A(n9), .B(n26), .Z(\ab[19][9] ) );
  NR2 U327 ( .A(n8), .B(n26), .Z(\ab[19][8] ) );
  NR2 U328 ( .A(n15), .B(n26), .Z(\ab[19][7] ) );
  NR2 U329 ( .A(n14), .B(n26), .Z(\ab[19][6] ) );
  NR2 U330 ( .A(n13), .B(n26), .Z(\ab[19][5] ) );
  NR2 U331 ( .A(n4), .B(n26), .Z(\ab[19][4] ) );
  NR2 U332 ( .A(n5), .B(n26), .Z(\ab[19][3] ) );
  NR2 U333 ( .A(n6), .B(n26), .Z(\ab[19][2] ) );
  NR2 U334 ( .A(n7), .B(n26), .Z(\ab[19][1] ) );
  NR2 U335 ( .A(n11), .B(n26), .Z(\ab[19][11] ) );
  NR2 U336 ( .A(n10), .B(n26), .Z(\ab[19][10] ) );
  NR2 U337 ( .A(n12), .B(n26), .Z(\ab[19][0] ) );
  NR2 U338 ( .A(n9), .B(n27), .Z(\ab[18][9] ) );
  NR2 U339 ( .A(n8), .B(n27), .Z(\ab[18][8] ) );
  NR2 U340 ( .A(n15), .B(n27), .Z(\ab[18][7] ) );
  NR2 U341 ( .A(n14), .B(n27), .Z(\ab[18][6] ) );
  NR2 U342 ( .A(n13), .B(n27), .Z(\ab[18][5] ) );
  NR2 U343 ( .A(n4), .B(n27), .Z(\ab[18][4] ) );
  NR2 U344 ( .A(n5), .B(n27), .Z(\ab[18][3] ) );
  NR2 U345 ( .A(n6), .B(n27), .Z(\ab[18][2] ) );
  NR2 U346 ( .A(n7), .B(n27), .Z(\ab[18][1] ) );
  NR2 U347 ( .A(n11), .B(n27), .Z(\ab[18][11] ) );
  NR2 U348 ( .A(n10), .B(n27), .Z(\ab[18][10] ) );
  NR2 U349 ( .A(n12), .B(n27), .Z(\ab[18][0] ) );
  NR2 U350 ( .A(n9), .B(n28), .Z(\ab[17][9] ) );
  NR2 U351 ( .A(n8), .B(n28), .Z(\ab[17][8] ) );
  NR2 U352 ( .A(n15), .B(n28), .Z(\ab[17][7] ) );
  NR2 U353 ( .A(n14), .B(n28), .Z(\ab[17][6] ) );
  NR2 U354 ( .A(n13), .B(n28), .Z(\ab[17][5] ) );
  NR2 U355 ( .A(n4), .B(n28), .Z(\ab[17][4] ) );
  NR2 U356 ( .A(n5), .B(n28), .Z(\ab[17][3] ) );
  NR2 U357 ( .A(n6), .B(n28), .Z(\ab[17][2] ) );
  NR2 U358 ( .A(n7), .B(n28), .Z(\ab[17][1] ) );
  NR2 U359 ( .A(n11), .B(n28), .Z(\ab[17][11] ) );
  NR2 U360 ( .A(n10), .B(n28), .Z(\ab[17][10] ) );
  NR2 U361 ( .A(n12), .B(n28), .Z(\ab[17][0] ) );
  NR2 U362 ( .A(n9), .B(n29), .Z(\ab[16][9] ) );
  NR2 U363 ( .A(n8), .B(n29), .Z(\ab[16][8] ) );
  NR2 U364 ( .A(n15), .B(n29), .Z(\ab[16][7] ) );
  NR2 U365 ( .A(n14), .B(n29), .Z(\ab[16][6] ) );
  NR2 U366 ( .A(n13), .B(n29), .Z(\ab[16][5] ) );
  NR2 U367 ( .A(n4), .B(n29), .Z(\ab[16][4] ) );
  NR2 U368 ( .A(n5), .B(n29), .Z(\ab[16][3] ) );
  NR2 U369 ( .A(n6), .B(n29), .Z(\ab[16][2] ) );
  NR2 U370 ( .A(n7), .B(n29), .Z(\ab[16][1] ) );
  NR2 U371 ( .A(n11), .B(n29), .Z(\ab[16][11] ) );
  NR2 U372 ( .A(n10), .B(n29), .Z(\ab[16][10] ) );
  NR2 U373 ( .A(n12), .B(n29), .Z(\ab[16][0] ) );
  NR2 U374 ( .A(n9), .B(n30), .Z(\ab[15][9] ) );
  NR2 U375 ( .A(n8), .B(n30), .Z(\ab[15][8] ) );
  NR2 U376 ( .A(n15), .B(n30), .Z(\ab[15][7] ) );
  NR2 U377 ( .A(n14), .B(n30), .Z(\ab[15][6] ) );
  NR2 U378 ( .A(n13), .B(n30), .Z(\ab[15][5] ) );
  NR2 U379 ( .A(n4), .B(n30), .Z(\ab[15][4] ) );
  NR2 U380 ( .A(n5), .B(n30), .Z(\ab[15][3] ) );
  NR2 U381 ( .A(n6), .B(n30), .Z(\ab[15][2] ) );
  NR2 U382 ( .A(n7), .B(n30), .Z(\ab[15][1] ) );
  NR2 U383 ( .A(n11), .B(n30), .Z(\ab[15][11] ) );
  NR2 U384 ( .A(n10), .B(n30), .Z(\ab[15][10] ) );
  NR2 U385 ( .A(n12), .B(n30), .Z(\ab[15][0] ) );
  NR2 U386 ( .A(n9), .B(n31), .Z(\ab[14][9] ) );
  NR2 U387 ( .A(n8), .B(n31), .Z(\ab[14][8] ) );
  NR2 U388 ( .A(n15), .B(n31), .Z(\ab[14][7] ) );
  NR2 U389 ( .A(n14), .B(n31), .Z(\ab[14][6] ) );
  NR2 U390 ( .A(n13), .B(n31), .Z(\ab[14][5] ) );
  NR2 U391 ( .A(n4), .B(n31), .Z(\ab[14][4] ) );
  NR2 U392 ( .A(n5), .B(n31), .Z(\ab[14][3] ) );
  NR2 U393 ( .A(n6), .B(n31), .Z(\ab[14][2] ) );
  NR2 U394 ( .A(n7), .B(n31), .Z(\ab[14][1] ) );
  NR2 U395 ( .A(n11), .B(n31), .Z(\ab[14][11] ) );
  NR2 U396 ( .A(n10), .B(n31), .Z(\ab[14][10] ) );
  NR2 U397 ( .A(n12), .B(n31), .Z(\ab[14][0] ) );
  NR2 U398 ( .A(n9), .B(n32), .Z(\ab[13][9] ) );
  NR2 U399 ( .A(n8), .B(n32), .Z(\ab[13][8] ) );
  NR2 U400 ( .A(n15), .B(n32), .Z(\ab[13][7] ) );
  NR2 U401 ( .A(n14), .B(n32), .Z(\ab[13][6] ) );
  NR2 U402 ( .A(n13), .B(n32), .Z(\ab[13][5] ) );
  NR2 U403 ( .A(n4), .B(n32), .Z(\ab[13][4] ) );
  NR2 U404 ( .A(n5), .B(n32), .Z(\ab[13][3] ) );
  NR2 U405 ( .A(n6), .B(n32), .Z(\ab[13][2] ) );
  NR2 U406 ( .A(n7), .B(n32), .Z(\ab[13][1] ) );
  NR2 U407 ( .A(n11), .B(n32), .Z(\ab[13][11] ) );
  NR2 U408 ( .A(n10), .B(n32), .Z(\ab[13][10] ) );
  NR2 U409 ( .A(n12), .B(n32), .Z(\ab[13][0] ) );
  NR2 U410 ( .A(n9), .B(n33), .Z(\ab[12][9] ) );
  NR2 U411 ( .A(n8), .B(n33), .Z(\ab[12][8] ) );
  NR2 U412 ( .A(n15), .B(n33), .Z(\ab[12][7] ) );
  NR2 U413 ( .A(n14), .B(n33), .Z(\ab[12][6] ) );
  NR2 U414 ( .A(n13), .B(n33), .Z(\ab[12][5] ) );
  NR2 U415 ( .A(n4), .B(n33), .Z(\ab[12][4] ) );
  NR2 U416 ( .A(n5), .B(n33), .Z(\ab[12][3] ) );
  NR2 U417 ( .A(n6), .B(n33), .Z(\ab[12][2] ) );
  NR2 U418 ( .A(n7), .B(n33), .Z(\ab[12][1] ) );
  NR2 U419 ( .A(n11), .B(n33), .Z(\ab[12][11] ) );
  NR2 U420 ( .A(n10), .B(n33), .Z(\ab[12][10] ) );
  NR2 U421 ( .A(n12), .B(n33), .Z(\ab[12][0] ) );
  NR2 U422 ( .A(n9), .B(n34), .Z(\ab[11][9] ) );
  NR2 U423 ( .A(n8), .B(n34), .Z(\ab[11][8] ) );
  NR2 U424 ( .A(n15), .B(n34), .Z(\ab[11][7] ) );
  NR2 U425 ( .A(n14), .B(n34), .Z(\ab[11][6] ) );
  NR2 U426 ( .A(n13), .B(n34), .Z(\ab[11][5] ) );
  NR2 U427 ( .A(n4), .B(n34), .Z(\ab[11][4] ) );
  NR2 U428 ( .A(n5), .B(n34), .Z(\ab[11][3] ) );
  NR2 U429 ( .A(n6), .B(n34), .Z(\ab[11][2] ) );
  NR2 U430 ( .A(n7), .B(n34), .Z(\ab[11][1] ) );
  NR2 U431 ( .A(n11), .B(n34), .Z(\ab[11][11] ) );
  NR2 U432 ( .A(n10), .B(n34), .Z(\ab[11][10] ) );
  NR2 U433 ( .A(n12), .B(n34), .Z(\ab[11][0] ) );
  NR2 U434 ( .A(n9), .B(n35), .Z(\ab[10][9] ) );
  NR2 U435 ( .A(n8), .B(n35), .Z(\ab[10][8] ) );
  NR2 U436 ( .A(n15), .B(n35), .Z(\ab[10][7] ) );
  NR2 U437 ( .A(n14), .B(n35), .Z(\ab[10][6] ) );
  NR2 U438 ( .A(n13), .B(n35), .Z(\ab[10][5] ) );
  NR2 U439 ( .A(n4), .B(n35), .Z(\ab[10][4] ) );
  NR2 U440 ( .A(n5), .B(n35), .Z(\ab[10][3] ) );
  NR2 U441 ( .A(n6), .B(n35), .Z(\ab[10][2] ) );
  NR2 U442 ( .A(n7), .B(n35), .Z(\ab[10][1] ) );
  NR2 U443 ( .A(n11), .B(n35), .Z(\ab[10][11] ) );
  NR2 U444 ( .A(n10), .B(n35), .Z(\ab[10][10] ) );
  NR2 U445 ( .A(n12), .B(n35), .Z(\ab[10][0] ) );
  NR2 U446 ( .A(n9), .B(n45), .Z(\ab[0][9] ) );
  NR2 U447 ( .A(n8), .B(n45), .Z(\ab[0][8] ) );
  NR2 U448 ( .A(n15), .B(n45), .Z(\ab[0][7] ) );
  NR2 U449 ( .A(n14), .B(n45), .Z(\ab[0][6] ) );
  NR2 U450 ( .A(n13), .B(n45), .Z(\ab[0][5] ) );
  NR2 U451 ( .A(n4), .B(n45), .Z(\ab[0][4] ) );
  NR2 U452 ( .A(n5), .B(n45), .Z(\ab[0][3] ) );
  NR2 U453 ( .A(n6), .B(n45), .Z(\ab[0][2] ) );
  NR2 U454 ( .A(n11), .B(n45), .Z(\ab[0][11] ) );
  NR2 U455 ( .A(n10), .B(n45), .Z(\ab[0][10] ) );
  AN3 U456 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U457 ( .A(n44), .B(n7), .Z(\ab[1][1] ) );
endmodule


module Poly_sqrt ( clock, reset, Datain, DataOut );
  input [30:0] Datain;
  output [16:0] DataOut;
  input clock, reset;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N70, N71, N72, N73, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425;
  tri   clock;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25;
  assign N36 = Datain[30];

  Poly_sqrt_DW01_add_0 add_1186 ( .A({1'b0, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19}), .B({1'b0, N39, N40, N41, N42, N43, N44, 
        N45, N46, N47, N48, N49, N50, N51}), .CI(1'b0), .SUM({N65, N64, N63, 
        N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52}) );
  Poly_sqrt_DW02_mult_0 mult_1183 ( .A({N36, Datain[29:0]}), .B({n20, n18, n19, 
        N10, N11, N12, N13, N14, N15, N16, N17, N18}), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25}) );
  FDS2L \DataOut_reg[16]  ( .CR(1'b1), .D(N73), .LD(n425), .CP(clock), .Q(
        DataOut[16]) );
  FDS2L \DataOut_reg[15]  ( .CR(1'b1), .D(N72), .LD(n425), .CP(clock), .Q(
        DataOut[15]) );
  FDS2L \DataOut_reg[14]  ( .CR(1'b1), .D(N71), .LD(n425), .CP(clock), .Q(
        DataOut[14]) );
  FDS2L \DataOut_reg[13]  ( .CR(1'b1), .D(N70), .LD(n425), .CP(clock), .Q(
        DataOut[13]) );
  FDS2L \DataOut_reg[12]  ( .CR(1'b1), .D(N64), .LD(n425), .CP(clock), .Q(
        DataOut[12]) );
  FDS2L \DataOut_reg[11]  ( .CR(1'b1), .D(N63), .LD(n425), .CP(clock), .Q(
        DataOut[11]) );
  FDS2L \DataOut_reg[10]  ( .CR(1'b1), .D(N62), .LD(n425), .CP(clock), .Q(
        DataOut[10]) );
  FDS2L \DataOut_reg[9]  ( .CR(1'b1), .D(N61), .LD(n425), .CP(clock), .Q(
        DataOut[9]) );
  FDS2L \DataOut_reg[8]  ( .CR(1'b1), .D(N60), .LD(n425), .CP(clock), .Q(
        DataOut[8]) );
  FDS2L \DataOut_reg[7]  ( .CR(1'b1), .D(N59), .LD(n425), .CP(clock), .Q(
        DataOut[7]) );
  FDS2L \DataOut_reg[6]  ( .CR(1'b1), .D(N58), .LD(n425), .CP(clock), .Q(
        DataOut[6]) );
  FDS2L \DataOut_reg[5]  ( .CR(1'b1), .D(N57), .LD(n425), .CP(clock), .Q(
        DataOut[5]) );
  FDS2L \DataOut_reg[4]  ( .CR(1'b1), .D(N56), .LD(n425), .CP(clock), .Q(
        DataOut[4]) );
  FDS2L \DataOut_reg[3]  ( .CR(1'b1), .D(N55), .LD(n425), .CP(clock), .Q(
        DataOut[3]) );
  FDS2L \DataOut_reg[2]  ( .CR(1'b1), .D(N54), .LD(n425), .CP(clock), .Q(
        DataOut[2]) );
  FDS2L \DataOut_reg[1]  ( .CR(1'b1), .D(N53), .LD(n425), .CP(clock), .Q(
        DataOut[1]) );
  FDS2L \DataOut_reg[0]  ( .CR(1'b1), .D(N52), .LD(n425), .CP(clock), .Q(
        DataOut[0]) );
  NR2 U20 ( .A(Datain[29]), .B(n26), .Z(n397) );
  AN4P U21 ( .A(n28), .B(n411), .C(n410), .D(n409), .Z(n18) );
  AN4P U22 ( .A(n127), .B(n411), .C(n410), .D(n409), .Z(n19) );
  AN4P U23 ( .A(n126), .B(n411), .C(n410), .D(n409), .Z(n20) );
  AN2P U24 ( .A(n323), .B(n322), .Z(n21) );
  AN2P U25 ( .A(n334), .B(Datain[27]), .Z(n22) );
  AN2P U26 ( .A(n407), .B(n406), .Z(n23) );
  OR2P U27 ( .A(Datain[26]), .B(Datain[27]), .Z(n24) );
  AN2P U28 ( .A(n342), .B(n341), .Z(n25) );
  ND2 U29 ( .A(n407), .B(n406), .Z(n127) );
  ND4 U30 ( .A(n394), .B(n393), .C(n392), .D(n391), .Z(N39) );
  ND3 U31 ( .A(n406), .B(n405), .C(n407), .Z(n136) );
  ND2 U32 ( .A(n406), .B(n405), .Z(n220) );
  ND2 U33 ( .A(n407), .B(n405), .Z(n290) );
  ND2 U34 ( .A(n407), .B(n406), .Z(n223) );
  ND2 U35 ( .A(n407), .B(n406), .Z(n252) );
  ND2 U36 ( .A(n406), .B(n405), .Z(n202) );
  ND2 U37 ( .A(n406), .B(n405), .Z(n203) );
  ND3 U38 ( .A(n406), .B(n405), .C(n407), .Z(n35) );
  ND2 U39 ( .A(n407), .B(n406), .Z(n30) );
  IVP U40 ( .A(Datain[27]), .Z(n407) );
  IVP U41 ( .A(Datain[26]), .Z(n406) );
  IVP U42 ( .A(Datain[25]), .Z(n405) );
  ND3 U43 ( .A(n347), .B(n346), .C(n345), .Z(N10) );
  ND2 U44 ( .A(n128), .B(n411), .Z(n347) );
  ND2 U45 ( .A(Datain[28]), .B(n411), .Z(n346) );
  ND2 U46 ( .A(n404), .B(n411), .Z(N11) );
  MUX21L U47 ( .A(n403), .B(n402), .S(Datain[28]), .Z(n404) );
  NR2 U48 ( .A(Datain[29]), .B(n21), .Z(n403) );
  ND4 U49 ( .A(n401), .B(n400), .C(n399), .D(n398), .Z(N12) );
  MUX21L U50 ( .A(n396), .B(n395), .S(Datain[29]), .Z(n401) );
  MUX21L U51 ( .A(N36), .B(n397), .S(Datain[28]), .Z(n400) );
  ND4 U52 ( .A(n369), .B(n368), .C(n367), .D(n366), .Z(N13) );
  MUX21L U53 ( .A(n360), .B(n361), .S(N36), .Z(n369) );
  MUX21L U54 ( .A(n362), .B(n363), .S(Datain[29]), .Z(n368) );
  MUX21L U55 ( .A(Datain[25]), .B(n406), .S(Datain[27]), .Z(n143) );
  ND2 U56 ( .A(n407), .B(n406), .Z(n138) );
  NR3 U57 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n126) );
  MUX21L U58 ( .A(n407), .B(Datain[26]), .S(Datain[25]), .Z(n150) );
  MUX21L U59 ( .A(n406), .B(n220), .S(Datain[27]), .Z(n146) );
  MUX21L U60 ( .A(n300), .B(Datain[25]), .S(Datain[26]), .Z(n157) );
  ND2 U61 ( .A(n219), .B(n218), .Z(n153) );
  MUX21L U62 ( .A(n230), .B(n407), .S(Datain[25]), .Z(n160) );
  MUX21L U63 ( .A(n281), .B(n280), .S(Datain[26]), .Z(n163) );
  IVP U64 ( .A(N36), .Z(n411) );
  IVP U65 ( .A(Datain[28]), .Z(n409) );
  IVP U66 ( .A(Datain[29]), .Z(n410) );
  NR3 U67 ( .A(N36), .B(Datain[28]), .C(n22), .Z(n355) );
  EO U68 ( .A(Datain[25]), .B(Datain[26]), .Z(n334) );
  NR3 U69 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n137) );
  NR3 U70 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n156) );
  NR3 U71 ( .A(Datain[29]), .B(n23), .C(N36), .Z(n372) );
  NR3 U72 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n106) );
  ND4 U73 ( .A(n359), .B(n358), .C(n357), .D(n356), .Z(N18) );
  MUX21L U74 ( .A(n350), .B(n351), .S(Datain[28]), .Z(n359) );
  MUX21L U75 ( .A(n352), .B(n353), .S(Datain[29]), .Z(n358) );
  MUX21L U76 ( .A(n355), .B(n354), .S(Datain[29]), .Z(n357) );
  AO7 U77 ( .A(Datain[25]), .B(Datain[26]), .C(Datain[27]), .Z(n139) );
  AO6 U78 ( .A(Datain[26]), .B(n407), .C(n217), .Z(n219) );
  NR2 U79 ( .A(Datain[25]), .B(Datain[27]), .Z(n217) );
  AO7 U80 ( .A(Datain[26]), .B(n405), .C(n407), .Z(n162) );
  AO7 U81 ( .A(Datain[27]), .B(n405), .C(n406), .Z(n151) );
  AO7 U82 ( .A(Datain[27]), .B(n406), .C(n207), .Z(n121) );
  ND2 U83 ( .A(Datain[25]), .B(Datain[26]), .Z(n207) );
  AO7 U84 ( .A(Datain[27]), .B(n405), .C(n406), .Z(n124) );
  AO7 U85 ( .A(Datain[25]), .B(Datain[26]), .C(n407), .Z(n123) );
  AO7 U86 ( .A(Datain[25]), .B(Datain[27]), .C(Datain[26]), .Z(n118) );
  AO7 U87 ( .A(Datain[25]), .B(Datain[27]), .C(Datain[26]), .Z(n89) );
  AO7 U88 ( .A(Datain[26]), .B(n407), .C(n405), .Z(n95) );
  AO7 U89 ( .A(Datain[25]), .B(n406), .C(Datain[27]), .Z(n76) );
  AO4 U90 ( .A(Datain[25]), .B(Datain[27]), .C(Datain[25]), .D(Datain[26]), 
        .Z(n79) );
  AO7 U91 ( .A(Datain[26]), .B(n407), .C(n337), .Z(n80) );
  ND2 U92 ( .A(Datain[25]), .B(Datain[27]), .Z(n337) );
  AO7 U93 ( .A(Datain[26]), .B(Datain[27]), .C(n405), .Z(n71) );
  AO7 U94 ( .A(Datain[25]), .B(n406), .C(n407), .Z(n73) );
  AO7 U95 ( .A(Datain[26]), .B(Datain[27]), .C(n405), .Z(n56) );
  AO7 U96 ( .A(Datain[25]), .B(Datain[27]), .C(n406), .Z(n49) );
  AO7 U97 ( .A(Datain[25]), .B(Datain[26]), .C(Datain[27]), .Z(n39) );
  AO7 U98 ( .A(Datain[25]), .B(Datain[26]), .C(n407), .Z(n42) );
  NR2 U99 ( .A(Datain[26]), .B(Datain[27]), .Z(n319) );
  NR2 U100 ( .A(Datain[25]), .B(Datain[26]), .Z(n321) );
  NR2 U101 ( .A(Datain[25]), .B(n406), .Z(n320) );
  NR2 U102 ( .A(Datain[26]), .B(Datain[27]), .Z(n291) );
  NR2 U103 ( .A(Datain[29]), .B(n287), .Z(n402) );
  EO U104 ( .A(Datain[26]), .B(Datain[27]), .Z(n26) );
  NR2 U105 ( .A(Datain[28]), .B(n408), .Z(n395) );
  IVP U106 ( .A(n130), .Z(n408) );
  AO7 U107 ( .A(Datain[25]), .B(Datain[26]), .C(Datain[27]), .Z(n130) );
  NR2 U108 ( .A(Datain[28]), .B(n318), .Z(n396) );
  ND3 U109 ( .A(Datain[27]), .B(n406), .C(Datain[25]), .Z(n318) );
  NR2 U110 ( .A(Datain[29]), .B(n24), .Z(n361) );
  NR2 U111 ( .A(Datain[27]), .B(n406), .Z(n158) );
  NR2 U112 ( .A(Datain[25]), .B(n406), .Z(n339) );
  NR2 U113 ( .A(Datain[25]), .B(n407), .Z(n340) );
  NR2 U114 ( .A(Datain[27]), .B(n405), .Z(n338) );
  NR2 U115 ( .A(Datain[26]), .B(Datain[27]), .Z(n304) );
  NR2 U116 ( .A(Datain[27]), .B(Datain[26]), .Z(n224) );
  NR2 U117 ( .A(Datain[25]), .B(n406), .Z(n226) );
  NR2 U118 ( .A(Datain[26]), .B(Datain[27]), .Z(n285) );
  NR2 U119 ( .A(Datain[26]), .B(n407), .Z(n286) );
  NR2 U120 ( .A(Datain[25]), .B(n406), .Z(n98) );
  ND2 U121 ( .A(n374), .B(n373), .Z(N38) );
  MUX21L U122 ( .A(n371), .B(n370), .S(N36), .Z(n374) );
  MUX21L U123 ( .A(n372), .B(Datain[29]), .S(Datain[28]), .Z(n373) );
  ND2 U124 ( .A(n349), .B(n348), .Z(N37) );
  ND2 U125 ( .A(Datain[28]), .B(n411), .Z(n349) );
  ND2 U126 ( .A(Datain[29]), .B(n411), .Z(n348) );
  MUX21L U127 ( .A(n405), .B(Datain[26]), .S(Datain[27]), .Z(n125) );
  MUX21L U128 ( .A(Datain[27]), .B(n221), .S(Datain[26]), .Z(n122) );
  MUX21L U129 ( .A(n183), .B(n405), .S(Datain[26]), .Z(n120) );
  ND4 U130 ( .A(n170), .B(Datain[29]), .C(n411), .D(n409), .Z(n356) );
  MUX21L U131 ( .A(Datain[25]), .B(n406), .S(Datain[27]), .Z(n170) );
  ND4 U132 ( .A(n61), .B(N36), .C(Datain[29]), .D(n409), .Z(n381) );
  AO7 U133 ( .A(Datain[25]), .B(n407), .C(Datain[26]), .Z(n61) );
  ND4 U134 ( .A(n32), .B(N36), .C(Datain[29]), .D(n409), .Z(n391) );
  NR2 U135 ( .A(Datain[26]), .B(Datain[27]), .Z(n32) );
  AN3 U136 ( .A(n169), .B(n411), .C(Datain[28]), .Z(n354) );
  AO7 U137 ( .A(Datain[25]), .B(Datain[27]), .C(Datain[26]), .Z(n169) );
  AN3 U138 ( .A(n166), .B(Datain[28]), .C(N36), .Z(n353) );
  ND2 U139 ( .A(n173), .B(n172), .Z(n166) );
  ND2 U140 ( .A(n407), .B(n406), .Z(n172) );
  EN U141 ( .A(Datain[25]), .B(Datain[26]), .Z(n173) );
  AN3 U142 ( .A(n171), .B(n411), .C(Datain[28]), .Z(n352) );
  ND2 U143 ( .A(n297), .B(n296), .Z(n171) );
  ND2 U144 ( .A(n407), .B(n405), .Z(n297) );
  ND2 U145 ( .A(Datain[26]), .B(n407), .Z(n296) );
  AN3 U146 ( .A(n167), .B(n410), .C(N36), .Z(n351) );
  ND2 U147 ( .A(n215), .B(n214), .Z(n167) );
  ND2 U148 ( .A(Datain[25]), .B(n406), .Z(n215) );
  ND2 U149 ( .A(Datain[27]), .B(n406), .Z(n214) );
  AN3 U150 ( .A(n168), .B(n410), .C(N36), .Z(n350) );
  ND2 U151 ( .A(n244), .B(n243), .Z(n168) );
  ND2 U152 ( .A(Datain[26]), .B(n407), .Z(n244) );
  ND2 U153 ( .A(Datain[26]), .B(n405), .Z(n243) );
  AN3 U154 ( .A(n131), .B(N36), .C(Datain[28]), .Z(n363) );
  ND3 U155 ( .A(n406), .B(n405), .C(n407), .Z(n131) );
  AN3 U156 ( .A(n134), .B(n411), .C(Datain[28]), .Z(n362) );
  AO7 U157 ( .A(Datain[25]), .B(Datain[27]), .C(n406), .Z(n134) );
  AN3 U158 ( .A(n133), .B(n409), .C(Datain[29]), .Z(n360) );
  ND2 U159 ( .A(n293), .B(n292), .Z(n133) );
  MUX21L U160 ( .A(n291), .B(Datain[27]), .S(Datain[25]), .Z(n293) );
  ND2 U161 ( .A(Datain[26]), .B(Datain[27]), .Z(n292) );
  EO U162 ( .A(Datain[25]), .B(Datain[26]), .Z(n141) );
  EO U163 ( .A(Datain[26]), .B(Datain[27]), .Z(n165) );
  EN U164 ( .A(Datain[25]), .B(Datain[27]), .Z(n154) );
  EO U165 ( .A(Datain[25]), .B(Datain[26]), .Z(n152) );
  ND2 U166 ( .A(n407), .B(n406), .Z(n29) );
  EO U167 ( .A(Datain[25]), .B(Datain[27]), .Z(n311) );
  EO U168 ( .A(Datain[26]), .B(Datain[27]), .Z(n238) );
  AN3 U169 ( .A(n62), .B(n410), .C(N36), .Z(n376) );
  ND2 U170 ( .A(Datain[27]), .B(n234), .Z(n62) );
  ND2 U171 ( .A(Datain[25]), .B(Datain[26]), .Z(n234) );
  AN3 U172 ( .A(n64), .B(n411), .C(Datain[29]), .Z(n375) );
  AO7 U173 ( .A(Datain[25]), .B(Datain[27]), .C(n406), .Z(n64) );
  EN U174 ( .A(Datain[25]), .B(Datain[26]), .Z(n91) );
  EO U175 ( .A(Datain[25]), .B(Datain[27]), .Z(n66) );
  EO U176 ( .A(Datain[25]), .B(Datain[27]), .Z(n54) );
  EO U177 ( .A(Datain[25]), .B(Datain[27]), .Z(n51) );
  MUX21L U178 ( .A(n290), .B(n407), .S(Datain[26]), .Z(n117) );
  MUX21L U179 ( .A(n223), .B(n222), .S(Datain[25]), .Z(n107) );
  MUX21L U180 ( .A(Datain[27]), .B(n282), .S(Datain[26]), .Z(n110) );
  MUX21L U181 ( .A(n336), .B(n407), .S(Datain[25]), .Z(n104) );
  MUX21L U182 ( .A(n252), .B(n251), .S(Datain[25]), .Z(n100) );
  MUX21L U183 ( .A(Datain[25]), .B(n406), .S(Datain[27]), .Z(n93) );
  ND2 U184 ( .A(n330), .B(n329), .Z(n96) );
  MUX21L U185 ( .A(n405), .B(n202), .S(Datain[27]), .Z(n82) );
  ND2 U186 ( .A(n407), .B(n405), .Z(n88) );
  MUX21L U187 ( .A(n406), .B(n203), .S(Datain[27]), .Z(n74) );
  ND2 U188 ( .A(n238), .B(n237), .Z(n75) );
  MUX21L U189 ( .A(Datain[26]), .B(Datain[27]), .S(Datain[25]), .Z(n72) );
  ND2 U190 ( .A(Datain[26]), .B(Datain[27]), .Z(n69) );
  ND4 U191 ( .A(n384), .B(n383), .C(n382), .D(n381), .Z(N43) );
  MUX21L U192 ( .A(n375), .B(n376), .S(Datain[28]), .Z(n384) );
  MUX21L U193 ( .A(Datain[26]), .B(n407), .S(Datain[25]), .Z(n52) );
  MUX21L U194 ( .A(Datain[27]), .B(n213), .S(Datain[26]), .Z(n40) );
  ND3 U195 ( .A(n135), .B(n409), .C(n410), .Z(n366) );
  MUX21L U196 ( .A(n407), .B(Datain[26]), .S(Datain[25]), .Z(n135) );
  ND3 U197 ( .A(n328), .B(n327), .C(n326), .Z(n119) );
  ND2 U198 ( .A(Datain[27]), .B(n405), .Z(n328) );
  ND2 U199 ( .A(n406), .B(n405), .Z(n327) );
  ND2 U200 ( .A(Datain[27]), .B(n406), .Z(n326) );
  ND3 U201 ( .A(Datain[26]), .B(n407), .C(Datain[25]), .Z(n77) );
  ND2 U202 ( .A(n325), .B(n324), .Z(n128) );
  ND2 U203 ( .A(n407), .B(n405), .Z(n325) );
  ND2 U204 ( .A(Datain[26]), .B(n407), .Z(n324) );
  ND2 U205 ( .A(Datain[29]), .B(n411), .Z(n345) );
  ND2 U206 ( .A(n129), .B(N36), .Z(n398) );
  NR3 U207 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n129) );
  ND2 U208 ( .A(N36), .B(n410), .Z(n399) );
  ND2 U209 ( .A(n315), .B(Datain[25]), .Z(n142) );
  EO U210 ( .A(Datain[26]), .B(Datain[27]), .Z(n315) );
  ND2 U211 ( .A(n265), .B(n264), .Z(n140) );
  ND2 U212 ( .A(Datain[25]), .B(n407), .Z(n265) );
  ND2 U213 ( .A(Datain[26]), .B(n407), .Z(n264) );
  ND2 U214 ( .A(Datain[25]), .B(Datain[27]), .Z(n280) );
  ND2 U215 ( .A(Datain[25]), .B(n407), .Z(n281) );
  ND2 U216 ( .A(Datain[26]), .B(n407), .Z(n230) );
  ND2 U217 ( .A(Datain[25]), .B(n407), .Z(n300) );
  ND2 U218 ( .A(Datain[27]), .B(n253), .Z(n161) );
  ND2 U219 ( .A(Datain[25]), .B(Datain[26]), .Z(n253) );
  ND2 U220 ( .A(n193), .B(n192), .Z(n159) );
  MUX21L U221 ( .A(n191), .B(n405), .S(Datain[27]), .Z(n193) );
  ND2 U222 ( .A(Datain[26]), .B(Datain[27]), .Z(n192) );
  NR2 U223 ( .A(Datain[26]), .B(n405), .Z(n191) );
  ND2 U224 ( .A(n299), .B(n298), .Z(n164) );
  ND2 U225 ( .A(Datain[25]), .B(n407), .Z(n298) );
  EN U226 ( .A(Datain[26]), .B(Datain[27]), .Z(n299) );
  ND2 U227 ( .A(n175), .B(n174), .Z(n144) );
  ND2 U228 ( .A(Datain[25]), .B(n407), .Z(n174) );
  EN U229 ( .A(Datain[26]), .B(Datain[27]), .Z(n175) );
  ND2 U230 ( .A(n247), .B(n246), .Z(n147) );
  MUX21L U231 ( .A(n406), .B(n245), .S(Datain[27]), .Z(n247) );
  ND2 U232 ( .A(Datain[25]), .B(n406), .Z(n246) );
  NR2 U233 ( .A(Datain[25]), .B(n406), .Z(n245) );
  ND2 U234 ( .A(n302), .B(n301), .Z(n149) );
  ND2 U235 ( .A(Datain[27]), .B(n405), .Z(n301) );
  EN U236 ( .A(Datain[26]), .B(Datain[27]), .Z(n302) );
  ND2 U237 ( .A(n198), .B(n197), .Z(n145) );
  MUX21L U238 ( .A(n196), .B(n407), .S(Datain[25]), .Z(n198) );
  ND2 U239 ( .A(Datain[26]), .B(n407), .Z(n197) );
  NR2 U240 ( .A(Datain[26]), .B(n407), .Z(n196) );
  ND2 U241 ( .A(n263), .B(n262), .Z(n148) );
  MUX21L U242 ( .A(Datain[25]), .B(n261), .S(Datain[26]), .Z(n263) );
  ND2 U243 ( .A(Datain[27]), .B(n406), .Z(n262) );
  NR2 U244 ( .A(Datain[25]), .B(Datain[27]), .Z(n261) );
  ND2 U245 ( .A(n260), .B(n259), .Z(n155) );
  ND2 U246 ( .A(n407), .B(n406), .Z(n259) );
  EN U247 ( .A(Datain[25]), .B(Datain[27]), .Z(n260) );
  ND2 U248 ( .A(Datain[26]), .B(Datain[27]), .Z(n316) );
  ND2 U249 ( .A(Datain[25]), .B(Datain[27]), .Z(n317) );
  ND2 U250 ( .A(Datain[27]), .B(n405), .Z(n183) );
  ND2 U251 ( .A(Datain[27]), .B(n405), .Z(n221) );
  ND2 U252 ( .A(Datain[25]), .B(Datain[27]), .Z(n282) );
  ND2 U253 ( .A(Datain[26]), .B(n407), .Z(n222) );
  ND2 U254 ( .A(Datain[27]), .B(n406), .Z(n251) );
  ND2 U255 ( .A(Datain[26]), .B(n407), .Z(n336) );
  ND2 U256 ( .A(Datain[25]), .B(n406), .Z(n329) );
  ND2 U257 ( .A(Datain[25]), .B(n407), .Z(n330) );
  ND2 U258 ( .A(Datain[27]), .B(n405), .Z(n237) );
  ND2 U259 ( .A(Datain[25]), .B(Datain[27]), .Z(n213) );
  ND2 U260 ( .A(n236), .B(n235), .Z(n114) );
  ND2 U261 ( .A(n407), .B(n405), .Z(n235) );
  EO U262 ( .A(Datain[26]), .B(Datain[27]), .Z(n236) );
  ND2 U263 ( .A(n201), .B(n200), .Z(n113) );
  MUX21L U264 ( .A(n199), .B(n405), .S(Datain[26]), .Z(n201) );
  ND2 U265 ( .A(Datain[27]), .B(n405), .Z(n200) );
  NR2 U266 ( .A(Datain[27]), .B(n405), .Z(n199) );
  ND2 U267 ( .A(n250), .B(n249), .Z(n115) );
  MUX21L U268 ( .A(Datain[25]), .B(n248), .S(Datain[26]), .Z(n250) );
  ND2 U269 ( .A(Datain[27]), .B(n406), .Z(n249) );
  NR2 U270 ( .A(Datain[25]), .B(Datain[27]), .Z(n248) );
  ND2 U271 ( .A(n272), .B(n271), .Z(n109) );
  MUX21L U272 ( .A(n270), .B(Datain[27]), .S(Datain[26]), .Z(n271) );
  AO2 U273 ( .A(Datain[25]), .B(Datain[27]), .C(Datain[25]), .D(Datain[26]), 
        .Z(n272) );
  NR2 U274 ( .A(Datain[25]), .B(Datain[27]), .Z(n270) );
  ND2 U275 ( .A(n258), .B(n257), .Z(n108) );
  EO U276 ( .A(Datain[25]), .B(Datain[27]), .Z(n258) );
  EO U277 ( .A(Datain[26]), .B(Datain[27]), .Z(n257) );
  ND2 U278 ( .A(n306), .B(n305), .Z(n111) );
  MUX21L U279 ( .A(Datain[25]), .B(n303), .S(Datain[26]), .Z(n305) );
  AO6 U280 ( .A(Datain[25]), .B(n407), .C(n304), .Z(n306) );
  NR2 U281 ( .A(Datain[25]), .B(n407), .Z(n303) );
  ND2 U282 ( .A(n186), .B(n185), .Z(n105) );
  MUX21L U283 ( .A(n406), .B(n184), .S(Datain[27]), .Z(n186) );
  ND2 U284 ( .A(n406), .B(n405), .Z(n185) );
  ND2 U285 ( .A(n335), .B(Datain[26]), .Z(n112) );
  EO U286 ( .A(Datain[25]), .B(Datain[27]), .Z(n335) );
  ND2 U287 ( .A(n269), .B(n268), .Z(n101) );
  MUX21L U288 ( .A(n405), .B(n267), .S(Datain[27]), .Z(n269) );
  ND2 U289 ( .A(n406), .B(n405), .Z(n268) );
  ND2 U290 ( .A(n228), .B(n227), .Z(n99) );
  MUX21L U291 ( .A(n225), .B(n226), .S(Datain[27]), .Z(n228) );
  ND2 U292 ( .A(n224), .B(n405), .Z(n227) );
  ND2 U293 ( .A(n284), .B(n283), .Z(n102) );
  ND2 U294 ( .A(Datain[26]), .B(Datain[25]), .Z(n284) );
  ND2 U295 ( .A(Datain[25]), .B(Datain[27]), .Z(n283) );
  ND2 U296 ( .A(n276), .B(n275), .Z(n94) );
  ND2 U297 ( .A(Datain[26]), .B(n405), .Z(n276) );
  ND2 U298 ( .A(Datain[27]), .B(n405), .Z(n275) );
  ND2 U299 ( .A(n210), .B(n209), .Z(n90) );
  MUX21L U300 ( .A(n406), .B(n208), .S(Datain[27]), .Z(n210) );
  ND2 U301 ( .A(n406), .B(n405), .Z(n209) );
  ND2 U302 ( .A(n255), .B(n254), .Z(n92) );
  ND2 U303 ( .A(n407), .B(n406), .Z(n254) );
  EO U304 ( .A(Datain[25]), .B(Datain[26]), .Z(n255) );
  ND2 U305 ( .A(n177), .B(n176), .Z(n81) );
  ND2 U306 ( .A(Datain[27]), .B(n406), .Z(n177) );
  ND2 U307 ( .A(Datain[27]), .B(n405), .Z(n176) );
  ND2 U308 ( .A(n273), .B(n406), .Z(n85) );
  EO U309 ( .A(Datain[25]), .B(Datain[27]), .Z(n273) );
  ND2 U310 ( .A(n232), .B(n231), .Z(n83) );
  ND2 U311 ( .A(Datain[27]), .B(n406), .Z(n231) );
  EO U312 ( .A(Datain[25]), .B(Datain[26]), .Z(n232) );
  ND2 U313 ( .A(n308), .B(n307), .Z(n87) );
  ND2 U314 ( .A(n407), .B(n406), .Z(n307) );
  EN U315 ( .A(Datain[25]), .B(Datain[27]), .Z(n308) );
  ND2 U316 ( .A(Datain[26]), .B(n405), .Z(n86) );
  ND2 U317 ( .A(n256), .B(Datain[25]), .Z(n84) );
  EO U318 ( .A(Datain[26]), .B(Datain[27]), .Z(n256) );
  ND2 U319 ( .A(n277), .B(Datain[25]), .Z(n78) );
  EN U320 ( .A(Datain[26]), .B(Datain[27]), .Z(n277) );
  ND2 U321 ( .A(n233), .B(Datain[26]), .Z(n68) );
  EO U322 ( .A(Datain[25]), .B(Datain[27]), .Z(n233) );
  ND2 U323 ( .A(n212), .B(n211), .Z(n67) );
  ND2 U324 ( .A(Datain[27]), .B(n406), .Z(n211) );
  EO U325 ( .A(Datain[25]), .B(Datain[27]), .Z(n212) );
  ND2 U326 ( .A(n274), .B(n407), .Z(n70) );
  EO U327 ( .A(Datain[25]), .B(Datain[26]), .Z(n274) );
  ND2 U328 ( .A(n310), .B(n309), .Z(n58) );
  ND2 U329 ( .A(Datain[27]), .B(n406), .Z(n310) );
  ND2 U330 ( .A(Datain[27]), .B(n405), .Z(n309) );
  ND2 U331 ( .A(n182), .B(n181), .Z(n53) );
  ND2 U332 ( .A(n407), .B(n406), .Z(n181) );
  EN U333 ( .A(Datain[25]), .B(Datain[27]), .Z(n182) );
  ND2 U334 ( .A(n279), .B(n278), .Z(n57) );
  ND2 U335 ( .A(n407), .B(n406), .Z(n278) );
  EN U336 ( .A(Datain[25]), .B(Datain[27]), .Z(n279) );
  ND2 U337 ( .A(Datain[25]), .B(n239), .Z(n55) );
  ND2 U338 ( .A(Datain[26]), .B(Datain[27]), .Z(n239) );
  ND2 U339 ( .A(n333), .B(n332), .Z(n59) );
  MUX21L U340 ( .A(n331), .B(n407), .S(Datain[25]), .Z(n333) );
  ND2 U341 ( .A(Datain[26]), .B(n407), .Z(n332) );
  NR2 U342 ( .A(Datain[26]), .B(n407), .Z(n331) );
  ND2 U343 ( .A(n190), .B(n189), .Z(n46) );
  MUX21L U344 ( .A(n188), .B(n407), .S(Datain[26]), .Z(n190) );
  ND2 U345 ( .A(Datain[25]), .B(Datain[26]), .Z(n189) );
  NR2 U346 ( .A(Datain[25]), .B(n407), .Z(n188) );
  ND2 U347 ( .A(n206), .B(n205), .Z(n47) );
  MUX21L U348 ( .A(n406), .B(n204), .S(Datain[27]), .Z(n206) );
  ND2 U349 ( .A(Datain[25]), .B(n406), .Z(n205) );
  NR2 U350 ( .A(Datain[25]), .B(n406), .Z(n204) );
  ND2 U351 ( .A(n289), .B(n288), .Z(n50) );
  MUX21L U352 ( .A(n286), .B(n287), .S(Datain[25]), .Z(n289) );
  ND2 U353 ( .A(n285), .B(Datain[25]), .Z(n288) );
  ND2 U354 ( .A(n314), .B(n313), .Z(n44) );
  MUX21L U355 ( .A(n312), .B(n407), .S(Datain[26]), .Z(n314) );
  ND2 U356 ( .A(Datain[25]), .B(Datain[26]), .Z(n313) );
  NR2 U357 ( .A(Datain[25]), .B(n407), .Z(n312) );
  ND2 U358 ( .A(n295), .B(n294), .Z(n43) );
  ND2 U359 ( .A(Datain[25]), .B(Datain[27]), .Z(n294) );
  EO U360 ( .A(Datain[26]), .B(Datain[27]), .Z(n295) );
  ND2 U361 ( .A(n242), .B(n241), .Z(n41) );
  MUX21L U362 ( .A(n240), .B(Datain[27]), .S(Datain[25]), .Z(n242) );
  ND2 U363 ( .A(Datain[26]), .B(Datain[27]), .Z(n241) );
  NR2 U364 ( .A(Datain[26]), .B(Datain[27]), .Z(n240) );
  ND2 U365 ( .A(n344), .B(n343), .Z(n45) );
  EN U366 ( .A(Datain[25]), .B(Datain[27]), .Z(n344) );
  EO U367 ( .A(Datain[26]), .B(Datain[27]), .Z(n343) );
  MUX21L U368 ( .A(n320), .B(n321), .S(Datain[27]), .Z(n323) );
  ND2 U369 ( .A(n319), .B(Datain[25]), .Z(n322) );
  MUX21L U370 ( .A(n338), .B(Datain[27]), .S(Datain[26]), .Z(n341) );
  NR2 U371 ( .A(n340), .B(n339), .Z(n342) );
  MUX21H U372 ( .A(n405), .B(n407), .S(Datain[26]), .Z(n27) );
  AN3 U373 ( .A(n407), .B(n406), .C(Datain[25]), .Z(n28) );
  MUX21L U374 ( .A(n364), .B(n365), .S(N36), .Z(n367) );
  AN3 U375 ( .A(Datain[29]), .B(n132), .C(Datain[28]), .Z(n364) );
  NR2 U376 ( .A(Datain[28]), .B(Datain[29]), .Z(n365) );
  NR3 U377 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n132) );
  MUX21L U378 ( .A(n216), .B(n405), .S(Datain[26]), .Z(n218) );
  MUX21L U379 ( .A(Datain[26]), .B(n266), .S(Datain[25]), .Z(n116) );
  ND2 U380 ( .A(Datain[26]), .B(n407), .Z(n266) );
  MUX21L U381 ( .A(Datain[25]), .B(Datain[26]), .S(Datain[27]), .Z(n103) );
  MUX21L U382 ( .A(n187), .B(n405), .S(Datain[26]), .Z(n97) );
  ND2 U383 ( .A(Datain[27]), .B(n405), .Z(n187) );
  MUX21L U384 ( .A(n380), .B(n379), .S(Datain[29]), .Z(n382) );
  AN3 U385 ( .A(n63), .B(n411), .C(Datain[28]), .Z(n379) );
  NR3 U386 ( .A(N36), .B(Datain[28]), .C(n25), .Z(n380) );
  NR3 U387 ( .A(Datain[27]), .B(Datain[25]), .C(Datain[26]), .Z(n63) );
  MUX21L U388 ( .A(n377), .B(n378), .S(Datain[29]), .Z(n383) );
  AN3 U389 ( .A(n65), .B(n411), .C(Datain[28]), .Z(n377) );
  AN3 U390 ( .A(n60), .B(Datain[28]), .C(N36), .Z(n378) );
  ND2 U391 ( .A(n311), .B(Datain[26]), .Z(n65) );
  MUX21L U392 ( .A(Datain[26]), .B(n229), .S(Datain[25]), .Z(n48) );
  ND2 U393 ( .A(Datain[26]), .B(n407), .Z(n229) );
  MUX21L U394 ( .A(n390), .B(n389), .S(Datain[29]), .Z(n392) );
  AN3 U395 ( .A(n36), .B(n411), .C(Datain[28]), .Z(n389) );
  NR3 U396 ( .A(N36), .B(Datain[28]), .C(n27), .Z(n390) );
  ND3 U397 ( .A(n406), .B(n405), .C(n407), .Z(n36) );
  MUX21L U398 ( .A(n387), .B(n388), .S(Datain[29]), .Z(n393) );
  AN3 U399 ( .A(n38), .B(n411), .C(Datain[28]), .Z(n387) );
  AN3 U400 ( .A(n31), .B(Datain[28]), .C(N36), .Z(n388) );
  ND2 U401 ( .A(n317), .B(n316), .Z(n38) );
  MUX21L U402 ( .A(n385), .B(n386), .S(Datain[28]), .Z(n394) );
  AN3 U403 ( .A(n37), .B(n411), .C(Datain[29]), .Z(n385) );
  AN3 U404 ( .A(n35), .B(n410), .C(N36), .Z(n386) );
  NR2 U405 ( .A(Datain[26]), .B(Datain[27]), .Z(n37) );
  ND2 U406 ( .A(n180), .B(n179), .Z(n60) );
  MUX21L U407 ( .A(Datain[25]), .B(n178), .S(Datain[26]), .Z(n180) );
  ND2 U408 ( .A(Datain[27]), .B(n406), .Z(n179) );
  NR2 U409 ( .A(Datain[25]), .B(Datain[27]), .Z(n178) );
  ND2 U410 ( .A(n195), .B(n194), .Z(n31) );
  ND2 U411 ( .A(Datain[25]), .B(Datain[27]), .Z(n195) );
  ND2 U412 ( .A(Datain[26]), .B(Datain[27]), .Z(n194) );
  MUX81P U413 ( .D0(n45), .D1(Datain[27]), .D2(n43), .D3(n40), .D4(n44), .D5(
        n41), .D6(n42), .D7(n39), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(
        N40) );
  MUX81P U414 ( .D0(n52), .D1(Datain[26]), .D2(n50), .D3(n47), .D4(n51), .D5(
        n48), .D6(n49), .D7(n46), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(
        N41) );
  MUX81P U415 ( .D0(n59), .D1(Datain[25]), .D2(n57), .D3(n54), .D4(n58), .D5(
        n55), .D6(n56), .D7(n53), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(
        N42) );
  MUX81P U416 ( .D0(n73), .D1(n69), .D2(n71), .D3(n67), .D4(n72), .D5(n68), 
        .D6(n70), .D7(n66), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(N44)
         );
  MUX81P U417 ( .D0(n80), .D1(n76), .D2(n78), .D3(n74), .D4(n79), .D5(n75), 
        .D6(n77), .D7(Datain[27]), .A(N36), .B(Datain[29]), .C(Datain[28]), 
        .Z(N45) );
  MUX81P U418 ( .D0(n88), .D1(n84), .D2(n86), .D3(n82), .D4(n87), .D5(n83), 
        .D6(n85), .D7(n81), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(N46)
         );
  MUX81P U419 ( .D0(n96), .D1(n92), .D2(n94), .D3(n90), .D4(n95), .D5(n91), 
        .D6(n93), .D7(n89), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(N47)
         );
  MUX81P U420 ( .D0(n104), .D1(n100), .D2(n102), .D3(n98), .D4(n103), .D5(n99), 
        .D6(n101), .D7(n97), .A(N36), .B(Datain[29]), .C(Datain[28]), .Z(N48)
         );
  MUX81P U421 ( .D0(n112), .D1(n108), .D2(n110), .D3(n106), .D4(n111), .D5(
        n107), .D6(n109), .D7(n105), .A(N36), .B(Datain[29]), .C(Datain[28]), 
        .Z(N49) );
  MUX81P U422 ( .D0(n119), .D1(n115), .D2(n117), .D3(n113), .D4(n118), .D5(
        n114), .D6(n116), .D7(Datain[27]), .A(N36), .B(Datain[29]), .C(
        Datain[28]), .Z(N50) );
  MUX81P U423 ( .D0(n125), .D1(n123), .D2(n28), .D3(n121), .D4(Datain[26]), 
        .D5(n122), .D6(n124), .D7(n120), .A(N36), .B(Datain[29]), .C(
        Datain[28]), .Z(N51) );
  MUX81P U424 ( .D0(n143), .D1(n139), .D2(n141), .D3(n137), .D4(n142), .D5(
        n138), .D6(n140), .D7(n136), .A(N36), .B(Datain[29]), .C(Datain[28]), 
        .Z(N14) );
  MUX81P U425 ( .D0(n150), .D1(n147), .D2(Datain[25]), .D3(n145), .D4(n149), 
        .D5(n146), .D6(n148), .D7(n144), .A(N36), .B(Datain[29]), .C(
        Datain[28]), .Z(N15) );
  MUX81P U426 ( .D0(n158), .D1(n154), .D2(n156), .D3(n152), .D4(n157), .D5(
        n153), .D6(n155), .D7(n151), .A(N36), .B(Datain[29]), .C(Datain[28]), 
        .Z(N16) );
  MUX81P U427 ( .D0(n165), .D1(n161), .D2(n163), .D3(Datain[25]), .D4(n164), 
        .D5(n160), .D6(n162), .D7(n159), .A(N36), .B(Datain[29]), .C(
        Datain[28]), .Z(N17) );
  AN2P U428 ( .A(Datain[25]), .B(Datain[26]), .Z(n184) );
  AN2P U429 ( .A(Datain[25]), .B(Datain[26]), .Z(n208) );
  AN2P U430 ( .A(Datain[25]), .B(Datain[27]), .Z(n216) );
  AN2P U431 ( .A(Datain[25]), .B(Datain[26]), .Z(n225) );
  AN2P U432 ( .A(Datain[25]), .B(Datain[26]), .Z(n267) );
  AN2P U433 ( .A(Datain[26]), .B(Datain[27]), .Z(n287) );
  AN2P U434 ( .A(n29), .B(Datain[29]), .Z(n370) );
  AN2P U435 ( .A(n30), .B(Datain[29]), .Z(n371) );
  IV U436 ( .A(reset), .Z(n425) );
  EN U437 ( .A(n412), .B(N35), .Z(N73) );
  AO5 U438 ( .A(N34), .B(n413), .C(N36), .Z(n412) );
  AO2 U439 ( .A(n414), .B(n415), .C(n416), .D(n417), .Z(n413) );
  IV U440 ( .A(N37), .Z(n415) );
  ND2 U441 ( .A(N33), .B(n418), .Z(n414) );
  EO U442 ( .A(n419), .B(n420), .Z(N72) );
  EN U443 ( .A(N34), .B(N36), .Z(n420) );
  AO4 U444 ( .A(N33), .B(n418), .C(N37), .D(n421), .Z(n419) );
  NR2 U445 ( .A(n416), .B(n417), .Z(n421) );
  IV U446 ( .A(n416), .Z(n418) );
  EO U447 ( .A(n422), .B(n416), .Z(N71) );
  AO2 U448 ( .A(N32), .B(N38), .C(n423), .D(N65), .Z(n416) );
  OR2 U449 ( .A(N32), .B(N38), .Z(n423) );
  EO U450 ( .A(n417), .B(N37), .Z(n422) );
  IV U451 ( .A(N33), .Z(n417) );
  EO U452 ( .A(N32), .B(n424), .Z(N70) );
  EO U453 ( .A(N65), .B(N38), .Z(n424) );
endmodule


module top_module_DW01_add_0 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  IVP U2 ( .A(n67), .Z(n14) );
  IVP U3 ( .A(n59), .Z(n12) );
  IVP U4 ( .A(n51), .Z(n10) );
  IVP U5 ( .A(n43), .Z(n8) );
  IVP U6 ( .A(n35), .Z(n6) );
  IVP U7 ( .A(n27), .Z(n4) );
  IVP U8 ( .A(n63), .Z(n13) );
  IVP U9 ( .A(n55), .Z(n11) );
  IVP U10 ( .A(n47), .Z(n9) );
  IVP U11 ( .A(n39), .Z(n7) );
  IVP U12 ( .A(n31), .Z(n5) );
  IVP U13 ( .A(n23), .Z(n3) );
  IVP U14 ( .A(n18), .Z(n1) );
  IVP U15 ( .A(n69), .Z(n15) );
  ND2 U16 ( .A(A[14]), .B(B[14]), .Z(n70) );
  IVP U17 ( .A(n19), .Z(n2) );
  EO U18 ( .A(n16), .B(B[29]), .Z(SUM[29]) );
  AO7 U19 ( .A(n17), .B(n2), .C(n18), .Z(n16) );
  EO U20 ( .A(n19), .B(n20), .Z(SUM[28]) );
  NR2 U21 ( .A(n1), .B(n17), .Z(n20) );
  NR2 U22 ( .A(B[28]), .B(A[28]), .Z(n17) );
  ND2 U23 ( .A(B[28]), .B(A[28]), .Z(n18) );
  AO7 U24 ( .A(n21), .B(n22), .C(n23), .Z(n19) );
  EN U25 ( .A(n22), .B(n24), .Z(SUM[27]) );
  NR2 U26 ( .A(n3), .B(n21), .Z(n24) );
  NR2 U27 ( .A(B[27]), .B(A[27]), .Z(n21) );
  ND2 U28 ( .A(B[27]), .B(A[27]), .Z(n23) );
  AO6 U29 ( .A(n4), .B(n25), .C(n26), .Z(n22) );
  EO U30 ( .A(n25), .B(n28), .Z(SUM[26]) );
  NR2 U31 ( .A(n26), .B(n27), .Z(n28) );
  NR2 U32 ( .A(B[26]), .B(A[26]), .Z(n27) );
  AN2 U33 ( .A(B[26]), .B(A[26]), .Z(n26) );
  AO7 U34 ( .A(n29), .B(n30), .C(n31), .Z(n25) );
  EN U35 ( .A(n30), .B(n32), .Z(SUM[25]) );
  NR2 U36 ( .A(n5), .B(n29), .Z(n32) );
  NR2 U37 ( .A(B[25]), .B(A[25]), .Z(n29) );
  ND2 U38 ( .A(B[25]), .B(A[25]), .Z(n31) );
  AO6 U39 ( .A(n6), .B(n33), .C(n34), .Z(n30) );
  EO U40 ( .A(n33), .B(n36), .Z(SUM[24]) );
  NR2 U41 ( .A(n34), .B(n35), .Z(n36) );
  NR2 U42 ( .A(B[24]), .B(A[24]), .Z(n35) );
  AN2 U43 ( .A(B[24]), .B(A[24]), .Z(n34) );
  AO7 U44 ( .A(n37), .B(n38), .C(n39), .Z(n33) );
  EN U45 ( .A(n38), .B(n40), .Z(SUM[23]) );
  NR2 U46 ( .A(n7), .B(n37), .Z(n40) );
  NR2 U47 ( .A(B[23]), .B(A[23]), .Z(n37) );
  ND2 U48 ( .A(B[23]), .B(A[23]), .Z(n39) );
  AO6 U49 ( .A(n8), .B(n41), .C(n42), .Z(n38) );
  EO U50 ( .A(n41), .B(n44), .Z(SUM[22]) );
  NR2 U51 ( .A(n42), .B(n43), .Z(n44) );
  NR2 U52 ( .A(B[22]), .B(A[22]), .Z(n43) );
  AN2 U53 ( .A(B[22]), .B(A[22]), .Z(n42) );
  AO7 U54 ( .A(n45), .B(n46), .C(n47), .Z(n41) );
  EN U55 ( .A(n46), .B(n48), .Z(SUM[21]) );
  NR2 U56 ( .A(n9), .B(n45), .Z(n48) );
  NR2 U57 ( .A(B[21]), .B(A[21]), .Z(n45) );
  ND2 U58 ( .A(B[21]), .B(A[21]), .Z(n47) );
  AO6 U59 ( .A(n10), .B(n49), .C(n50), .Z(n46) );
  EO U60 ( .A(n49), .B(n52), .Z(SUM[20]) );
  NR2 U61 ( .A(n50), .B(n51), .Z(n52) );
  NR2 U62 ( .A(B[20]), .B(A[20]), .Z(n51) );
  AN2 U63 ( .A(B[20]), .B(A[20]), .Z(n50) );
  AO7 U64 ( .A(n53), .B(n54), .C(n55), .Z(n49) );
  EN U65 ( .A(n54), .B(n56), .Z(SUM[19]) );
  NR2 U66 ( .A(n11), .B(n53), .Z(n56) );
  NR2 U67 ( .A(B[19]), .B(A[19]), .Z(n53) );
  ND2 U68 ( .A(B[19]), .B(A[19]), .Z(n55) );
  AO6 U69 ( .A(n12), .B(n57), .C(n58), .Z(n54) );
  EO U70 ( .A(n57), .B(n60), .Z(SUM[18]) );
  NR2 U71 ( .A(n58), .B(n59), .Z(n60) );
  NR2 U72 ( .A(B[18]), .B(A[18]), .Z(n59) );
  AN2 U73 ( .A(B[18]), .B(A[18]), .Z(n58) );
  AO7 U74 ( .A(n61), .B(n62), .C(n63), .Z(n57) );
  EN U75 ( .A(n62), .B(n64), .Z(SUM[17]) );
  NR2 U76 ( .A(n13), .B(n61), .Z(n64) );
  NR2 U77 ( .A(B[17]), .B(A[17]), .Z(n61) );
  ND2 U78 ( .A(B[17]), .B(A[17]), .Z(n63) );
  AO6 U79 ( .A(n14), .B(n65), .C(n66), .Z(n62) );
  EO U80 ( .A(n65), .B(n68), .Z(SUM[16]) );
  NR2 U81 ( .A(n66), .B(n67), .Z(n68) );
  NR2 U82 ( .A(B[16]), .B(A[16]), .Z(n67) );
  AN2 U83 ( .A(B[16]), .B(A[16]), .Z(n66) );
  AO7 U84 ( .A(n69), .B(n70), .C(n71), .Z(n65) );
  EO U85 ( .A(n72), .B(n70), .Z(SUM[15]) );
  ND2 U86 ( .A(n15), .B(n71), .Z(n72) );
  ND2 U87 ( .A(B[15]), .B(A[15]), .Z(n71) );
  NR2 U88 ( .A(B[15]), .B(A[15]), .Z(n69) );
endmodule


module top_module_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [14:0] A;
  input [16:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][16] ,
         \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] ,
         \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] ,
         \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] ,
         \ab[12][0] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][16] ,
         \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] ,
         \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] ,
         \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] ,
         \ab[7][0] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][16] ,
         \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] ,
         \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] ,
         \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[14][0] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] ,
         \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] ,
         \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] ,
         \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] ,
         \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] ,
         \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[29] , \A2[28] , \A2[27] , \A2[26] ,
         \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] ,
         \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  tri   [14:0] A;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  top_module_DW01_add_0 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \SUMB[14][0] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[29] , 
        \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , 
        \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , 
        \A2[14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[31:17], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S4_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\SUMB[14][0] ) );
  FA1A S4_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S5_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\ab[13][16] ), .CO(
        \CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S4_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S3_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\ab[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S4_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S4_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S3_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\ab[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S4_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S4_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S3_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\ab[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S4_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(
        \CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S4_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S3_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\ab[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S4_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S4_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(
        \CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S3_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\ab[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S4_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S4_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S3_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\ab[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S4_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(
        \CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S4_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(
        \CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S3_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\ab[6][16] ), .CO(
        \CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S3_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\ab[5][16] ), .CO(
        \CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S3_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\ab[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S3_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\ab[3][16] ), .CO(
        \CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S3_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\ab[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S3_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  EO U2 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A1[14] ) );
  EO U3 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A1[15] ) );
  EO U4 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A1[16] ) );
  EO U5 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A1[17] ) );
  EO U6 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A1[18] ) );
  EO U7 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A1[19] ) );
  EO U8 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A1[20] ) );
  EO U9 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A1[21] ) );
  EO U10 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A1[22] ) );
  EO U11 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A1[23] ) );
  EO U12 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A1[24] ) );
  EO U13 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A1[25] ) );
  EO U14 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A1[26] ) );
  EO U15 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A1[27] ) );
  EO U16 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A1[28] ) );
  EO U17 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A1[13] ) );
  EO U18 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U19 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U20 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U21 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U22 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U23 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U24 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U25 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U26 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U27 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U28 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U29 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U30 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U31 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  IVP U32 ( .A(B[8]), .Z(n11) );
  IVP U33 ( .A(B[7]), .Z(n12) );
  IVP U34 ( .A(B[6]), .Z(n13) );
  IVP U35 ( .A(B[5]), .Z(n14) );
  IVP U36 ( .A(B[4]), .Z(n15) );
  IVP U37 ( .A(B[3]), .Z(n16) );
  IVP U38 ( .A(B[2]), .Z(n17) );
  IVP U39 ( .A(B[10]), .Z(n9) );
  IVP U40 ( .A(B[9]), .Z(n10) );
  IVP U41 ( .A(B[12]), .Z(n7) );
  IVP U42 ( .A(B[11]), .Z(n8) );
  IVP U43 ( .A(B[14]), .Z(n5) );
  IVP U44 ( .A(B[13]), .Z(n6) );
  IVP U45 ( .A(B[16]), .Z(n3) );
  IVP U46 ( .A(B[15]), .Z(n4) );
  IVP U47 ( .A(B[1]), .Z(n18) );
  IVP U48 ( .A(B[0]), .Z(n19) );
  EO U49 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  AN2P U50 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A2[14] ) );
  AN2P U51 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A2[16] ) );
  AN2P U52 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A2[17] ) );
  AN2P U53 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A2[18] ) );
  AN2P U54 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A2[19] ) );
  AN2P U55 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A2[20] ) );
  AN2P U56 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A2[21] ) );
  AN2P U57 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A2[22] ) );
  AN2P U58 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A2[23] ) );
  AN2P U59 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A2[24] ) );
  AN2P U60 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A2[25] ) );
  AN2P U61 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A2[26] ) );
  AN2P U62 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A2[27] ) );
  AN2P U63 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A2[28] ) );
  AN2P U64 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A2[29] ) );
  AN2P U65 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U66 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U67 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U68 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U69 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U70 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U71 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U72 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U73 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U74 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U75 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U76 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U77 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U78 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U79 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U80 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A2[15] ) );
  NR2 U82 ( .A(n22), .B(n10), .Z(\ab[9][9] ) );
  NR2 U83 ( .A(n22), .B(n11), .Z(\ab[9][8] ) );
  NR2 U84 ( .A(n22), .B(n12), .Z(\ab[9][7] ) );
  NR2 U85 ( .A(n22), .B(n13), .Z(\ab[9][6] ) );
  NR2 U86 ( .A(n22), .B(n14), .Z(\ab[9][5] ) );
  NR2 U87 ( .A(n22), .B(n15), .Z(\ab[9][4] ) );
  NR2 U88 ( .A(n22), .B(n16), .Z(\ab[9][3] ) );
  NR2 U89 ( .A(n22), .B(n17), .Z(\ab[9][2] ) );
  NR2 U90 ( .A(n22), .B(n18), .Z(\ab[9][1] ) );
  NR2 U91 ( .A(n22), .B(n3), .Z(\ab[9][16] ) );
  NR2 U92 ( .A(n22), .B(n4), .Z(\ab[9][15] ) );
  NR2 U93 ( .A(n22), .B(n5), .Z(\ab[9][14] ) );
  NR2 U94 ( .A(n22), .B(n6), .Z(\ab[9][13] ) );
  NR2 U95 ( .A(n22), .B(n7), .Z(\ab[9][12] ) );
  NR2 U96 ( .A(n22), .B(n8), .Z(\ab[9][11] ) );
  NR2 U97 ( .A(n22), .B(n9), .Z(\ab[9][10] ) );
  NR2 U98 ( .A(n22), .B(n19), .Z(\ab[9][0] ) );
  IV U99 ( .A(A[9]), .Z(n22) );
  NR2 U100 ( .A(n10), .B(n23), .Z(\ab[8][9] ) );
  NR2 U101 ( .A(n11), .B(n23), .Z(\ab[8][8] ) );
  NR2 U102 ( .A(n12), .B(n23), .Z(\ab[8][7] ) );
  NR2 U103 ( .A(n13), .B(n23), .Z(\ab[8][6] ) );
  NR2 U104 ( .A(n14), .B(n23), .Z(\ab[8][5] ) );
  NR2 U105 ( .A(n15), .B(n23), .Z(\ab[8][4] ) );
  NR2 U106 ( .A(n16), .B(n23), .Z(\ab[8][3] ) );
  NR2 U107 ( .A(n17), .B(n23), .Z(\ab[8][2] ) );
  NR2 U108 ( .A(n18), .B(n23), .Z(\ab[8][1] ) );
  NR2 U109 ( .A(n3), .B(n23), .Z(\ab[8][16] ) );
  NR2 U110 ( .A(n4), .B(n23), .Z(\ab[8][15] ) );
  NR2 U111 ( .A(n5), .B(n23), .Z(\ab[8][14] ) );
  NR2 U112 ( .A(n6), .B(n23), .Z(\ab[8][13] ) );
  NR2 U113 ( .A(n7), .B(n23), .Z(\ab[8][12] ) );
  NR2 U114 ( .A(n8), .B(n23), .Z(\ab[8][11] ) );
  NR2 U115 ( .A(n9), .B(n23), .Z(\ab[8][10] ) );
  NR2 U116 ( .A(n19), .B(n23), .Z(\ab[8][0] ) );
  IV U117 ( .A(A[8]), .Z(n23) );
  NR2 U118 ( .A(n10), .B(n24), .Z(\ab[7][9] ) );
  NR2 U119 ( .A(n11), .B(n24), .Z(\ab[7][8] ) );
  NR2 U120 ( .A(n12), .B(n24), .Z(\ab[7][7] ) );
  NR2 U121 ( .A(n13), .B(n24), .Z(\ab[7][6] ) );
  NR2 U122 ( .A(n14), .B(n24), .Z(\ab[7][5] ) );
  NR2 U123 ( .A(n15), .B(n24), .Z(\ab[7][4] ) );
  NR2 U124 ( .A(n16), .B(n24), .Z(\ab[7][3] ) );
  NR2 U125 ( .A(n17), .B(n24), .Z(\ab[7][2] ) );
  NR2 U126 ( .A(n18), .B(n24), .Z(\ab[7][1] ) );
  NR2 U127 ( .A(n3), .B(n24), .Z(\ab[7][16] ) );
  NR2 U128 ( .A(n4), .B(n24), .Z(\ab[7][15] ) );
  NR2 U129 ( .A(n5), .B(n24), .Z(\ab[7][14] ) );
  NR2 U130 ( .A(n6), .B(n24), .Z(\ab[7][13] ) );
  NR2 U131 ( .A(n7), .B(n24), .Z(\ab[7][12] ) );
  NR2 U132 ( .A(n8), .B(n24), .Z(\ab[7][11] ) );
  NR2 U133 ( .A(n9), .B(n24), .Z(\ab[7][10] ) );
  NR2 U134 ( .A(n19), .B(n24), .Z(\ab[7][0] ) );
  IV U135 ( .A(A[7]), .Z(n24) );
  NR2 U136 ( .A(n10), .B(n25), .Z(\ab[6][9] ) );
  NR2 U137 ( .A(n11), .B(n25), .Z(\ab[6][8] ) );
  NR2 U138 ( .A(n12), .B(n25), .Z(\ab[6][7] ) );
  NR2 U139 ( .A(n13), .B(n25), .Z(\ab[6][6] ) );
  NR2 U140 ( .A(n14), .B(n25), .Z(\ab[6][5] ) );
  NR2 U141 ( .A(n15), .B(n25), .Z(\ab[6][4] ) );
  NR2 U142 ( .A(n16), .B(n25), .Z(\ab[6][3] ) );
  NR2 U143 ( .A(n17), .B(n25), .Z(\ab[6][2] ) );
  NR2 U144 ( .A(n18), .B(n25), .Z(\ab[6][1] ) );
  NR2 U145 ( .A(n3), .B(n25), .Z(\ab[6][16] ) );
  NR2 U146 ( .A(n4), .B(n25), .Z(\ab[6][15] ) );
  NR2 U147 ( .A(n5), .B(n25), .Z(\ab[6][14] ) );
  NR2 U148 ( .A(n6), .B(n25), .Z(\ab[6][13] ) );
  NR2 U149 ( .A(n7), .B(n25), .Z(\ab[6][12] ) );
  NR2 U150 ( .A(n8), .B(n25), .Z(\ab[6][11] ) );
  NR2 U151 ( .A(n9), .B(n25), .Z(\ab[6][10] ) );
  NR2 U152 ( .A(n19), .B(n25), .Z(\ab[6][0] ) );
  IV U153 ( .A(A[6]), .Z(n25) );
  NR2 U154 ( .A(n10), .B(n26), .Z(\ab[5][9] ) );
  NR2 U155 ( .A(n11), .B(n26), .Z(\ab[5][8] ) );
  NR2 U156 ( .A(n12), .B(n26), .Z(\ab[5][7] ) );
  NR2 U157 ( .A(n13), .B(n26), .Z(\ab[5][6] ) );
  NR2 U158 ( .A(n14), .B(n26), .Z(\ab[5][5] ) );
  NR2 U159 ( .A(n15), .B(n26), .Z(\ab[5][4] ) );
  NR2 U160 ( .A(n16), .B(n26), .Z(\ab[5][3] ) );
  NR2 U161 ( .A(n17), .B(n26), .Z(\ab[5][2] ) );
  NR2 U162 ( .A(n18), .B(n26), .Z(\ab[5][1] ) );
  NR2 U163 ( .A(n3), .B(n26), .Z(\ab[5][16] ) );
  NR2 U164 ( .A(n4), .B(n26), .Z(\ab[5][15] ) );
  NR2 U165 ( .A(n5), .B(n26), .Z(\ab[5][14] ) );
  NR2 U166 ( .A(n6), .B(n26), .Z(\ab[5][13] ) );
  NR2 U167 ( .A(n7), .B(n26), .Z(\ab[5][12] ) );
  NR2 U168 ( .A(n8), .B(n26), .Z(\ab[5][11] ) );
  NR2 U169 ( .A(n9), .B(n26), .Z(\ab[5][10] ) );
  NR2 U170 ( .A(n19), .B(n26), .Z(\ab[5][0] ) );
  IV U171 ( .A(A[5]), .Z(n26) );
  NR2 U172 ( .A(n10), .B(n27), .Z(\ab[4][9] ) );
  NR2 U173 ( .A(n11), .B(n27), .Z(\ab[4][8] ) );
  NR2 U174 ( .A(n12), .B(n27), .Z(\ab[4][7] ) );
  NR2 U175 ( .A(n13), .B(n27), .Z(\ab[4][6] ) );
  NR2 U176 ( .A(n14), .B(n27), .Z(\ab[4][5] ) );
  NR2 U177 ( .A(n15), .B(n27), .Z(\ab[4][4] ) );
  NR2 U178 ( .A(n16), .B(n27), .Z(\ab[4][3] ) );
  NR2 U179 ( .A(n17), .B(n27), .Z(\ab[4][2] ) );
  NR2 U180 ( .A(n18), .B(n27), .Z(\ab[4][1] ) );
  NR2 U181 ( .A(n3), .B(n27), .Z(\ab[4][16] ) );
  NR2 U182 ( .A(n4), .B(n27), .Z(\ab[4][15] ) );
  NR2 U183 ( .A(n5), .B(n27), .Z(\ab[4][14] ) );
  NR2 U184 ( .A(n6), .B(n27), .Z(\ab[4][13] ) );
  NR2 U185 ( .A(n7), .B(n27), .Z(\ab[4][12] ) );
  NR2 U186 ( .A(n8), .B(n27), .Z(\ab[4][11] ) );
  NR2 U187 ( .A(n9), .B(n27), .Z(\ab[4][10] ) );
  NR2 U188 ( .A(n19), .B(n27), .Z(\ab[4][0] ) );
  IV U189 ( .A(A[4]), .Z(n27) );
  NR2 U190 ( .A(n10), .B(n28), .Z(\ab[3][9] ) );
  NR2 U191 ( .A(n11), .B(n28), .Z(\ab[3][8] ) );
  NR2 U192 ( .A(n12), .B(n28), .Z(\ab[3][7] ) );
  NR2 U193 ( .A(n13), .B(n28), .Z(\ab[3][6] ) );
  NR2 U194 ( .A(n14), .B(n28), .Z(\ab[3][5] ) );
  NR2 U195 ( .A(n15), .B(n28), .Z(\ab[3][4] ) );
  NR2 U196 ( .A(n16), .B(n28), .Z(\ab[3][3] ) );
  NR2 U197 ( .A(n17), .B(n28), .Z(\ab[3][2] ) );
  NR2 U198 ( .A(n18), .B(n28), .Z(\ab[3][1] ) );
  NR2 U199 ( .A(n3), .B(n28), .Z(\ab[3][16] ) );
  NR2 U200 ( .A(n4), .B(n28), .Z(\ab[3][15] ) );
  NR2 U201 ( .A(n5), .B(n28), .Z(\ab[3][14] ) );
  NR2 U202 ( .A(n6), .B(n28), .Z(\ab[3][13] ) );
  NR2 U203 ( .A(n7), .B(n28), .Z(\ab[3][12] ) );
  NR2 U204 ( .A(n8), .B(n28), .Z(\ab[3][11] ) );
  NR2 U205 ( .A(n9), .B(n28), .Z(\ab[3][10] ) );
  NR2 U206 ( .A(n19), .B(n28), .Z(\ab[3][0] ) );
  IV U207 ( .A(A[3]), .Z(n28) );
  NR2 U208 ( .A(n10), .B(n29), .Z(\ab[2][9] ) );
  NR2 U209 ( .A(n11), .B(n29), .Z(\ab[2][8] ) );
  NR2 U210 ( .A(n12), .B(n29), .Z(\ab[2][7] ) );
  NR2 U211 ( .A(n13), .B(n29), .Z(\ab[2][6] ) );
  NR2 U212 ( .A(n14), .B(n29), .Z(\ab[2][5] ) );
  NR2 U213 ( .A(n15), .B(n29), .Z(\ab[2][4] ) );
  NR2 U214 ( .A(n16), .B(n29), .Z(\ab[2][3] ) );
  NR2 U215 ( .A(n17), .B(n29), .Z(\ab[2][2] ) );
  NR2 U216 ( .A(n18), .B(n29), .Z(\ab[2][1] ) );
  NR2 U217 ( .A(n3), .B(n29), .Z(\ab[2][16] ) );
  NR2 U218 ( .A(n4), .B(n29), .Z(\ab[2][15] ) );
  NR2 U219 ( .A(n5), .B(n29), .Z(\ab[2][14] ) );
  NR2 U220 ( .A(n6), .B(n29), .Z(\ab[2][13] ) );
  NR2 U221 ( .A(n7), .B(n29), .Z(\ab[2][12] ) );
  NR2 U222 ( .A(n8), .B(n29), .Z(\ab[2][11] ) );
  NR2 U223 ( .A(n9), .B(n29), .Z(\ab[2][10] ) );
  NR2 U224 ( .A(n19), .B(n29), .Z(\ab[2][0] ) );
  IV U225 ( .A(A[2]), .Z(n29) );
  NR2 U226 ( .A(n10), .B(n30), .Z(\ab[1][9] ) );
  NR2 U227 ( .A(n11), .B(n30), .Z(\ab[1][8] ) );
  NR2 U228 ( .A(n12), .B(n30), .Z(\ab[1][7] ) );
  NR2 U229 ( .A(n13), .B(n30), .Z(\ab[1][6] ) );
  NR2 U230 ( .A(n14), .B(n30), .Z(\ab[1][5] ) );
  NR2 U231 ( .A(n15), .B(n30), .Z(\ab[1][4] ) );
  NR2 U232 ( .A(n16), .B(n30), .Z(\ab[1][3] ) );
  NR2 U233 ( .A(n17), .B(n30), .Z(\ab[1][2] ) );
  NR2 U234 ( .A(n3), .B(n30), .Z(\ab[1][16] ) );
  NR2 U235 ( .A(n4), .B(n30), .Z(\ab[1][15] ) );
  NR2 U236 ( .A(n5), .B(n30), .Z(\ab[1][14] ) );
  NR2 U237 ( .A(n6), .B(n30), .Z(\ab[1][13] ) );
  NR2 U238 ( .A(n7), .B(n30), .Z(\ab[1][12] ) );
  NR2 U239 ( .A(n8), .B(n30), .Z(\ab[1][11] ) );
  NR2 U240 ( .A(n9), .B(n30), .Z(\ab[1][10] ) );
  NR2 U241 ( .A(n10), .B(n31), .Z(\ab[14][9] ) );
  NR2 U242 ( .A(n11), .B(n31), .Z(\ab[14][8] ) );
  NR2 U243 ( .A(n12), .B(n31), .Z(\ab[14][7] ) );
  NR2 U244 ( .A(n13), .B(n31), .Z(\ab[14][6] ) );
  NR2 U245 ( .A(n14), .B(n31), .Z(\ab[14][5] ) );
  NR2 U246 ( .A(n15), .B(n31), .Z(\ab[14][4] ) );
  NR2 U247 ( .A(n16), .B(n31), .Z(\ab[14][3] ) );
  NR2 U248 ( .A(n17), .B(n31), .Z(\ab[14][2] ) );
  NR2 U249 ( .A(n18), .B(n31), .Z(\ab[14][1] ) );
  NR2 U250 ( .A(n3), .B(n31), .Z(\ab[14][16] ) );
  NR2 U251 ( .A(n4), .B(n31), .Z(\ab[14][15] ) );
  NR2 U252 ( .A(n5), .B(n31), .Z(\ab[14][14] ) );
  NR2 U253 ( .A(n6), .B(n31), .Z(\ab[14][13] ) );
  NR2 U254 ( .A(n7), .B(n31), .Z(\ab[14][12] ) );
  NR2 U255 ( .A(n8), .B(n31), .Z(\ab[14][11] ) );
  NR2 U256 ( .A(n9), .B(n31), .Z(\ab[14][10] ) );
  NR2 U257 ( .A(n19), .B(n31), .Z(\ab[14][0] ) );
  IV U258 ( .A(A[14]), .Z(n31) );
  NR2 U259 ( .A(n10), .B(n32), .Z(\ab[13][9] ) );
  NR2 U260 ( .A(n11), .B(n32), .Z(\ab[13][8] ) );
  NR2 U261 ( .A(n12), .B(n32), .Z(\ab[13][7] ) );
  NR2 U262 ( .A(n13), .B(n32), .Z(\ab[13][6] ) );
  NR2 U263 ( .A(n14), .B(n32), .Z(\ab[13][5] ) );
  NR2 U264 ( .A(n15), .B(n32), .Z(\ab[13][4] ) );
  NR2 U265 ( .A(n16), .B(n32), .Z(\ab[13][3] ) );
  NR2 U266 ( .A(n17), .B(n32), .Z(\ab[13][2] ) );
  NR2 U267 ( .A(n18), .B(n32), .Z(\ab[13][1] ) );
  NR2 U268 ( .A(n3), .B(n32), .Z(\ab[13][16] ) );
  NR2 U269 ( .A(n4), .B(n32), .Z(\ab[13][15] ) );
  NR2 U270 ( .A(n5), .B(n32), .Z(\ab[13][14] ) );
  NR2 U271 ( .A(n6), .B(n32), .Z(\ab[13][13] ) );
  NR2 U272 ( .A(n7), .B(n32), .Z(\ab[13][12] ) );
  NR2 U273 ( .A(n8), .B(n32), .Z(\ab[13][11] ) );
  NR2 U274 ( .A(n9), .B(n32), .Z(\ab[13][10] ) );
  NR2 U275 ( .A(n19), .B(n32), .Z(\ab[13][0] ) );
  IV U276 ( .A(A[13]), .Z(n32) );
  NR2 U277 ( .A(n10), .B(n33), .Z(\ab[12][9] ) );
  NR2 U278 ( .A(n11), .B(n33), .Z(\ab[12][8] ) );
  NR2 U279 ( .A(n12), .B(n33), .Z(\ab[12][7] ) );
  NR2 U280 ( .A(n13), .B(n33), .Z(\ab[12][6] ) );
  NR2 U281 ( .A(n14), .B(n33), .Z(\ab[12][5] ) );
  NR2 U282 ( .A(n15), .B(n33), .Z(\ab[12][4] ) );
  NR2 U283 ( .A(n16), .B(n33), .Z(\ab[12][3] ) );
  NR2 U284 ( .A(n17), .B(n33), .Z(\ab[12][2] ) );
  NR2 U285 ( .A(n18), .B(n33), .Z(\ab[12][1] ) );
  NR2 U286 ( .A(n3), .B(n33), .Z(\ab[12][16] ) );
  NR2 U287 ( .A(n4), .B(n33), .Z(\ab[12][15] ) );
  NR2 U288 ( .A(n5), .B(n33), .Z(\ab[12][14] ) );
  NR2 U289 ( .A(n6), .B(n33), .Z(\ab[12][13] ) );
  NR2 U290 ( .A(n7), .B(n33), .Z(\ab[12][12] ) );
  NR2 U291 ( .A(n8), .B(n33), .Z(\ab[12][11] ) );
  NR2 U292 ( .A(n9), .B(n33), .Z(\ab[12][10] ) );
  NR2 U293 ( .A(n19), .B(n33), .Z(\ab[12][0] ) );
  IV U294 ( .A(A[12]), .Z(n33) );
  NR2 U295 ( .A(n10), .B(n34), .Z(\ab[11][9] ) );
  NR2 U296 ( .A(n11), .B(n34), .Z(\ab[11][8] ) );
  NR2 U297 ( .A(n12), .B(n34), .Z(\ab[11][7] ) );
  NR2 U298 ( .A(n13), .B(n34), .Z(\ab[11][6] ) );
  NR2 U299 ( .A(n14), .B(n34), .Z(\ab[11][5] ) );
  NR2 U300 ( .A(n15), .B(n34), .Z(\ab[11][4] ) );
  NR2 U301 ( .A(n16), .B(n34), .Z(\ab[11][3] ) );
  NR2 U302 ( .A(n17), .B(n34), .Z(\ab[11][2] ) );
  NR2 U303 ( .A(n18), .B(n34), .Z(\ab[11][1] ) );
  NR2 U304 ( .A(n3), .B(n34), .Z(\ab[11][16] ) );
  NR2 U305 ( .A(n4), .B(n34), .Z(\ab[11][15] ) );
  NR2 U306 ( .A(n5), .B(n34), .Z(\ab[11][14] ) );
  NR2 U307 ( .A(n6), .B(n34), .Z(\ab[11][13] ) );
  NR2 U308 ( .A(n7), .B(n34), .Z(\ab[11][12] ) );
  NR2 U309 ( .A(n8), .B(n34), .Z(\ab[11][11] ) );
  NR2 U310 ( .A(n9), .B(n34), .Z(\ab[11][10] ) );
  NR2 U311 ( .A(n19), .B(n34), .Z(\ab[11][0] ) );
  IV U312 ( .A(A[11]), .Z(n34) );
  NR2 U313 ( .A(n10), .B(n35), .Z(\ab[10][9] ) );
  NR2 U314 ( .A(n11), .B(n35), .Z(\ab[10][8] ) );
  NR2 U315 ( .A(n12), .B(n35), .Z(\ab[10][7] ) );
  NR2 U316 ( .A(n13), .B(n35), .Z(\ab[10][6] ) );
  NR2 U317 ( .A(n14), .B(n35), .Z(\ab[10][5] ) );
  NR2 U318 ( .A(n15), .B(n35), .Z(\ab[10][4] ) );
  NR2 U319 ( .A(n16), .B(n35), .Z(\ab[10][3] ) );
  NR2 U320 ( .A(n17), .B(n35), .Z(\ab[10][2] ) );
  NR2 U321 ( .A(n18), .B(n35), .Z(\ab[10][1] ) );
  NR2 U322 ( .A(n3), .B(n35), .Z(\ab[10][16] ) );
  NR2 U323 ( .A(n4), .B(n35), .Z(\ab[10][15] ) );
  NR2 U324 ( .A(n5), .B(n35), .Z(\ab[10][14] ) );
  NR2 U325 ( .A(n6), .B(n35), .Z(\ab[10][13] ) );
  NR2 U326 ( .A(n7), .B(n35), .Z(\ab[10][12] ) );
  NR2 U327 ( .A(n8), .B(n35), .Z(\ab[10][11] ) );
  NR2 U328 ( .A(n9), .B(n35), .Z(\ab[10][10] ) );
  NR2 U329 ( .A(n19), .B(n35), .Z(\ab[10][0] ) );
  IV U330 ( .A(A[10]), .Z(n35) );
  NR2 U331 ( .A(n10), .B(n36), .Z(\ab[0][9] ) );
  NR2 U332 ( .A(n11), .B(n36), .Z(\ab[0][8] ) );
  NR2 U333 ( .A(n12), .B(n36), .Z(\ab[0][7] ) );
  NR2 U334 ( .A(n13), .B(n36), .Z(\ab[0][6] ) );
  NR2 U335 ( .A(n14), .B(n36), .Z(\ab[0][5] ) );
  NR2 U336 ( .A(n15), .B(n36), .Z(\ab[0][4] ) );
  NR2 U337 ( .A(n16), .B(n36), .Z(\ab[0][3] ) );
  NR2 U338 ( .A(n17), .B(n36), .Z(\ab[0][2] ) );
  NR2 U339 ( .A(n3), .B(n36), .Z(\ab[0][16] ) );
  NR2 U340 ( .A(n4), .B(n36), .Z(\ab[0][15] ) );
  NR2 U341 ( .A(n5), .B(n36), .Z(\ab[0][14] ) );
  NR2 U342 ( .A(n6), .B(n36), .Z(\ab[0][13] ) );
  NR2 U343 ( .A(n7), .B(n36), .Z(\ab[0][12] ) );
  NR2 U344 ( .A(n8), .B(n36), .Z(\ab[0][11] ) );
  NR2 U345 ( .A(n9), .B(n36), .Z(\ab[0][10] ) );
  IV U346 ( .A(A[0]), .Z(n36) );
  AN3 U347 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U348 ( .A(n30), .B(n18), .Z(\ab[1][1] ) );
  IV U349 ( .A(A[1]), .Z(n30) );
endmodule


module top_module_DW01_add_1 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72;

  IVP U2 ( .A(n67), .Z(n14) );
  IVP U3 ( .A(n59), .Z(n12) );
  IVP U4 ( .A(n51), .Z(n10) );
  IVP U5 ( .A(n43), .Z(n8) );
  IVP U6 ( .A(n35), .Z(n6) );
  IVP U7 ( .A(n27), .Z(n4) );
  IVP U8 ( .A(n63), .Z(n13) );
  IVP U9 ( .A(n55), .Z(n11) );
  IVP U10 ( .A(n47), .Z(n9) );
  IVP U11 ( .A(n39), .Z(n7) );
  IVP U12 ( .A(n31), .Z(n5) );
  IVP U13 ( .A(n23), .Z(n3) );
  IVP U14 ( .A(n18), .Z(n1) );
  IVP U15 ( .A(n69), .Z(n15) );
  ND2 U16 ( .A(A[14]), .B(B[14]), .Z(n70) );
  IVP U17 ( .A(n19), .Z(n2) );
  EO U18 ( .A(n16), .B(B[29]), .Z(SUM[29]) );
  AO7 U19 ( .A(n17), .B(n2), .C(n18), .Z(n16) );
  EO U20 ( .A(n19), .B(n20), .Z(SUM[28]) );
  NR2 U21 ( .A(n1), .B(n17), .Z(n20) );
  NR2 U22 ( .A(B[28]), .B(A[28]), .Z(n17) );
  ND2 U23 ( .A(B[28]), .B(A[28]), .Z(n18) );
  AO7 U24 ( .A(n21), .B(n22), .C(n23), .Z(n19) );
  EN U25 ( .A(n22), .B(n24), .Z(SUM[27]) );
  NR2 U26 ( .A(n3), .B(n21), .Z(n24) );
  NR2 U27 ( .A(B[27]), .B(A[27]), .Z(n21) );
  ND2 U28 ( .A(B[27]), .B(A[27]), .Z(n23) );
  AO6 U29 ( .A(n4), .B(n25), .C(n26), .Z(n22) );
  EO U30 ( .A(n25), .B(n28), .Z(SUM[26]) );
  NR2 U31 ( .A(n26), .B(n27), .Z(n28) );
  NR2 U32 ( .A(B[26]), .B(A[26]), .Z(n27) );
  AN2 U33 ( .A(B[26]), .B(A[26]), .Z(n26) );
  AO7 U34 ( .A(n29), .B(n30), .C(n31), .Z(n25) );
  EN U35 ( .A(n30), .B(n32), .Z(SUM[25]) );
  NR2 U36 ( .A(n5), .B(n29), .Z(n32) );
  NR2 U37 ( .A(B[25]), .B(A[25]), .Z(n29) );
  ND2 U38 ( .A(B[25]), .B(A[25]), .Z(n31) );
  AO6 U39 ( .A(n6), .B(n33), .C(n34), .Z(n30) );
  EO U40 ( .A(n33), .B(n36), .Z(SUM[24]) );
  NR2 U41 ( .A(n34), .B(n35), .Z(n36) );
  NR2 U42 ( .A(B[24]), .B(A[24]), .Z(n35) );
  AN2 U43 ( .A(B[24]), .B(A[24]), .Z(n34) );
  AO7 U44 ( .A(n37), .B(n38), .C(n39), .Z(n33) );
  EN U45 ( .A(n38), .B(n40), .Z(SUM[23]) );
  NR2 U46 ( .A(n7), .B(n37), .Z(n40) );
  NR2 U47 ( .A(B[23]), .B(A[23]), .Z(n37) );
  ND2 U48 ( .A(B[23]), .B(A[23]), .Z(n39) );
  AO6 U49 ( .A(n8), .B(n41), .C(n42), .Z(n38) );
  EO U50 ( .A(n41), .B(n44), .Z(SUM[22]) );
  NR2 U51 ( .A(n42), .B(n43), .Z(n44) );
  NR2 U52 ( .A(B[22]), .B(A[22]), .Z(n43) );
  AN2 U53 ( .A(B[22]), .B(A[22]), .Z(n42) );
  AO7 U54 ( .A(n45), .B(n46), .C(n47), .Z(n41) );
  EN U55 ( .A(n46), .B(n48), .Z(SUM[21]) );
  NR2 U56 ( .A(n9), .B(n45), .Z(n48) );
  NR2 U57 ( .A(B[21]), .B(A[21]), .Z(n45) );
  ND2 U58 ( .A(B[21]), .B(A[21]), .Z(n47) );
  AO6 U59 ( .A(n10), .B(n49), .C(n50), .Z(n46) );
  EO U60 ( .A(n49), .B(n52), .Z(SUM[20]) );
  NR2 U61 ( .A(n50), .B(n51), .Z(n52) );
  NR2 U62 ( .A(B[20]), .B(A[20]), .Z(n51) );
  AN2 U63 ( .A(B[20]), .B(A[20]), .Z(n50) );
  AO7 U64 ( .A(n53), .B(n54), .C(n55), .Z(n49) );
  EN U65 ( .A(n54), .B(n56), .Z(SUM[19]) );
  NR2 U66 ( .A(n11), .B(n53), .Z(n56) );
  NR2 U67 ( .A(B[19]), .B(A[19]), .Z(n53) );
  ND2 U68 ( .A(B[19]), .B(A[19]), .Z(n55) );
  AO6 U69 ( .A(n12), .B(n57), .C(n58), .Z(n54) );
  EO U70 ( .A(n57), .B(n60), .Z(SUM[18]) );
  NR2 U71 ( .A(n58), .B(n59), .Z(n60) );
  NR2 U72 ( .A(B[18]), .B(A[18]), .Z(n59) );
  AN2 U73 ( .A(B[18]), .B(A[18]), .Z(n58) );
  AO7 U74 ( .A(n61), .B(n62), .C(n63), .Z(n57) );
  EN U75 ( .A(n62), .B(n64), .Z(SUM[17]) );
  NR2 U76 ( .A(n13), .B(n61), .Z(n64) );
  NR2 U77 ( .A(B[17]), .B(A[17]), .Z(n61) );
  ND2 U78 ( .A(B[17]), .B(A[17]), .Z(n63) );
  AO6 U79 ( .A(n14), .B(n65), .C(n66), .Z(n62) );
  EO U80 ( .A(n65), .B(n68), .Z(SUM[16]) );
  NR2 U81 ( .A(n66), .B(n67), .Z(n68) );
  NR2 U82 ( .A(B[16]), .B(A[16]), .Z(n67) );
  AN2 U83 ( .A(B[16]), .B(A[16]), .Z(n66) );
  AO7 U84 ( .A(n69), .B(n70), .C(n71), .Z(n65) );
  EO U85 ( .A(n72), .B(n70), .Z(SUM[15]) );
  ND2 U86 ( .A(n15), .B(n71), .Z(n72) );
  ND2 U87 ( .A(B[15]), .B(A[15]), .Z(n71) );
  NR2 U88 ( .A(B[15]), .B(A[15]), .Z(n69) );
endmodule


module top_module_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [14:0] A;
  input [16:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[14][16] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][16] ,
         \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] ,
         \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] ,
         \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] ,
         \ab[12][0] , \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] ,
         \ab[11][12] , \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] ,
         \ab[11][7] , \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] ,
         \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][16] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][16] ,
         \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] ,
         \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] ,
         \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] ,
         \ab[7][0] , \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] ,
         \ab[6][12] , \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] ,
         \ab[6][7] , \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] ,
         \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][16] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][16] ,
         \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] ,
         \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] ,
         \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] ,
         \ab[2][0] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] ,
         \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] ,
         \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] ,
         \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] ,
         \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[14][0] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] ,
         \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] ,
         \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] ,
         \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] ,
         \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] ,
         \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] ,
         \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][15] , \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] ,
         \SUMB[4][11] , \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] ,
         \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] ,
         \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][15] , \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] ,
         \SUMB[1][11] , \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] ,
         \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] ,
         \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[29] , \A2[28] , \A2[27] , \A2[26] ,
         \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] ,
         \A2[18] , \A2[17] , \A2[16] , \A2[15] , \A2[14] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36;
  tri   [14:0] A;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  top_module_DW01_add_1 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , 
        \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , 
        \SUMB[14][0] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , 
        \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[29] , 
        \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , 
        \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , 
        \A2[14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[31:17], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  FA1A S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA1A S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA1A S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA1A S4_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(
        \CARRYB[14][0] ), .S(\SUMB[14][0] ) );
  FA1A S4_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(
        \CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA1A S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA1A S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA1A S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA1A S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA1A S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA1A S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA1A S5_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\ab[13][16] ), .CO(
        \CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA1A S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA1A S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA1A S4_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA1A S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA1A S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA1A S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA1A S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA1A S3_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\ab[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA1A S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA1A S4_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA1A S4_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA1A S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA1A S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA1A S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA1A S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA1A S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA1A S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA1A S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA1A S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA1A S3_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\ab[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA1A S4_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA1A S4_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA1A S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA1A S3_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\ab[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA1A S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA1A S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA1A S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA1A S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA1A S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA1A S4_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(
        \CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA1A S4_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), .CO(
        \CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA1A S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA1A S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA1A S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA1A S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA1A S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA1A S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA1A S3_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\ab[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA1A S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA1A S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA1A S4_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA1A S4_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(
        \CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA1A S3_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\ab[8][16] ), .CO(
        \CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA1A S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA1A S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA1A S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA1A S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA1A S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA1A S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA1A S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA1A S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA1A S4_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(
        \CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA1A S4_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(
        \CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA1A S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA1A S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA1A S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA1A S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA1A S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA1A S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA1A S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA1A S3_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\ab[7][16] ), .CO(
        \CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA1A S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA1A S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA1A S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA1A S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA1A S4_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(
        \CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA1A S4_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(
        \CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA1A S3_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\ab[6][16] ), .CO(
        \CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA1A S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA1A S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA1A S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA1A S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA1A S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA1A S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA1A S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA1A S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA1A S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA1A S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA1A S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), .CO(
        \CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA1A S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA1A S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA1A S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA1A S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA1A S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA1A S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA1A S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA1A S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA1A S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA1A S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA1A S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA1A S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA1A S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA1A S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA1A S3_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\ab[5][16] ), .CO(
        \CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA1A S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA1A S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA1A S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA1A S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA1A S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA1A S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA1A S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA1A S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA1A S3_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\ab[4][16] ), .CO(
        \CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA1A S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA1A S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA1A S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA1A S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA1A S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA1A S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA1A S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA1A S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA1A S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA1A S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA1A S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA1A S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA1A S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA1A S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA1A S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA1A S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA1A S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA1A S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA1A S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA1A S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA1A S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA1A S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA1A S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA1A S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA1A S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA1A S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA1A S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA1A S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA1A S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA1A S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA1A S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA1A S3_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\ab[3][16] ), .CO(
        \CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA1A S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA1A S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA1A S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA1A S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA1A S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA1A S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA1A S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA1A S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA1A S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA1A S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA1A S3_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\ab[2][16] ), .CO(
        \CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA1A S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA1A S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA1A S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA1A S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA1A S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA1A S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA1A S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA1A S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA1A S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA1A S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA1A S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA1A S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA1A S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA1A S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA1A S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA1A S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA1A S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA1A S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA1A S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA1A S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA1A S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA1A S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA1A S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA1A S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA1A S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA1A S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA1A S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA1A S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA1A S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA1A S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA1A S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA1A S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA1A S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA1A S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA1A S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA1A S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA1A S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA1A S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA1A S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA1A S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA1A S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA1A S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA1A S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA1A S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA1A S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA1A S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA1A S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA1A S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA1A S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA1A S3_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\ab[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  EO U2 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A1[14] ) );
  EO U3 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A1[15] ) );
  EO U4 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A1[16] ) );
  EO U5 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A1[17] ) );
  EO U6 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A1[18] ) );
  EO U7 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A1[19] ) );
  EO U8 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A1[20] ) );
  EO U9 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A1[21] ) );
  EO U10 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A1[22] ) );
  EO U11 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A1[23] ) );
  EO U12 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A1[24] ) );
  EO U13 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A1[25] ) );
  EO U14 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A1[26] ) );
  EO U15 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A1[27] ) );
  EO U16 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A1[28] ) );
  EO U17 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A1[13] ) );
  EO U18 ( .A(\ab[0][16] ), .B(\ab[1][15] ), .Z(\SUMB[1][15] ) );
  EO U19 ( .A(\ab[0][15] ), .B(\ab[1][14] ), .Z(\SUMB[1][14] ) );
  EO U20 ( .A(\ab[0][14] ), .B(\ab[1][13] ), .Z(\SUMB[1][13] ) );
  EO U21 ( .A(\ab[0][13] ), .B(\ab[1][12] ), .Z(\SUMB[1][12] ) );
  EO U22 ( .A(\ab[0][12] ), .B(\ab[1][11] ), .Z(\SUMB[1][11] ) );
  EO U23 ( .A(\ab[0][11] ), .B(\ab[1][10] ), .Z(\SUMB[1][10] ) );
  EO U24 ( .A(\ab[0][10] ), .B(\ab[1][9] ), .Z(\SUMB[1][9] ) );
  EO U25 ( .A(\ab[0][9] ), .B(\ab[1][8] ), .Z(\SUMB[1][8] ) );
  EO U26 ( .A(\ab[0][8] ), .B(\ab[1][7] ), .Z(\SUMB[1][7] ) );
  EO U27 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Z(\SUMB[1][6] ) );
  EO U28 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Z(\SUMB[1][5] ) );
  EO U29 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Z(\SUMB[1][4] ) );
  EO U30 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Z(\SUMB[1][3] ) );
  EO U31 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  IVP U32 ( .A(B[8]), .Z(n11) );
  IVP U33 ( .A(B[7]), .Z(n12) );
  IVP U34 ( .A(B[6]), .Z(n13) );
  IVP U35 ( .A(B[5]), .Z(n14) );
  IVP U36 ( .A(B[4]), .Z(n15) );
  IVP U37 ( .A(B[3]), .Z(n16) );
  IVP U38 ( .A(B[2]), .Z(n17) );
  IVP U39 ( .A(B[10]), .Z(n9) );
  IVP U40 ( .A(B[9]), .Z(n10) );
  IVP U41 ( .A(B[12]), .Z(n7) );
  IVP U42 ( .A(B[11]), .Z(n8) );
  IVP U43 ( .A(B[14]), .Z(n5) );
  IVP U44 ( .A(B[13]), .Z(n6) );
  IVP U45 ( .A(B[16]), .Z(n3) );
  IVP U46 ( .A(B[15]), .Z(n4) );
  IVP U47 ( .A(B[1]), .Z(n18) );
  IVP U48 ( .A(B[0]), .Z(n19) );
  EO U49 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  AN2P U50 ( .A(\CARRYB[14][0] ), .B(\SUMB[14][1] ), .Z(\A2[14] ) );
  AN2P U51 ( .A(\CARRYB[14][2] ), .B(\SUMB[14][3] ), .Z(\A2[16] ) );
  AN2P U52 ( .A(\CARRYB[14][3] ), .B(\SUMB[14][4] ), .Z(\A2[17] ) );
  AN2P U53 ( .A(\CARRYB[14][4] ), .B(\SUMB[14][5] ), .Z(\A2[18] ) );
  AN2P U54 ( .A(\CARRYB[14][5] ), .B(\SUMB[14][6] ), .Z(\A2[19] ) );
  AN2P U55 ( .A(\CARRYB[14][6] ), .B(\SUMB[14][7] ), .Z(\A2[20] ) );
  AN2P U56 ( .A(\CARRYB[14][7] ), .B(\SUMB[14][8] ), .Z(\A2[21] ) );
  AN2P U57 ( .A(\CARRYB[14][8] ), .B(\SUMB[14][9] ), .Z(\A2[22] ) );
  AN2P U58 ( .A(\CARRYB[14][9] ), .B(\SUMB[14][10] ), .Z(\A2[23] ) );
  AN2P U59 ( .A(\CARRYB[14][10] ), .B(\SUMB[14][11] ), .Z(\A2[24] ) );
  AN2P U60 ( .A(\CARRYB[14][11] ), .B(\SUMB[14][12] ), .Z(\A2[25] ) );
  AN2P U61 ( .A(\CARRYB[14][12] ), .B(\SUMB[14][13] ), .Z(\A2[26] ) );
  AN2P U62 ( .A(\CARRYB[14][13] ), .B(\SUMB[14][14] ), .Z(\A2[27] ) );
  AN2P U63 ( .A(\CARRYB[14][14] ), .B(\SUMB[14][15] ), .Z(\A2[28] ) );
  AN2P U64 ( .A(\CARRYB[14][15] ), .B(\ab[14][16] ), .Z(\A2[29] ) );
  AN2P U65 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  AN2P U66 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  AN2P U67 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\CARRYB[1][3] ) );
  AN2P U68 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\CARRYB[1][4] ) );
  AN2P U69 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\CARRYB[1][5] ) );
  AN2P U70 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\CARRYB[1][6] ) );
  AN2P U71 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\CARRYB[1][7] ) );
  AN2P U72 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\CARRYB[1][8] ) );
  AN2P U73 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\CARRYB[1][9] ) );
  AN2P U74 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\CARRYB[1][10] ) );
  AN2P U75 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\CARRYB[1][11] ) );
  AN2P U76 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\CARRYB[1][12] ) );
  AN2P U77 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\CARRYB[1][13] ) );
  AN2P U78 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\CARRYB[1][14] ) );
  AN2P U79 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\CARRYB[1][15] ) );
  AN2P U80 ( .A(\CARRYB[14][1] ), .B(\SUMB[14][2] ), .Z(\A2[15] ) );
  NR2 U82 ( .A(n22), .B(n10), .Z(\ab[9][9] ) );
  NR2 U83 ( .A(n22), .B(n11), .Z(\ab[9][8] ) );
  NR2 U84 ( .A(n22), .B(n12), .Z(\ab[9][7] ) );
  NR2 U85 ( .A(n22), .B(n13), .Z(\ab[9][6] ) );
  NR2 U86 ( .A(n22), .B(n14), .Z(\ab[9][5] ) );
  NR2 U87 ( .A(n22), .B(n15), .Z(\ab[9][4] ) );
  NR2 U88 ( .A(n22), .B(n16), .Z(\ab[9][3] ) );
  NR2 U89 ( .A(n22), .B(n17), .Z(\ab[9][2] ) );
  NR2 U90 ( .A(n22), .B(n18), .Z(\ab[9][1] ) );
  NR2 U91 ( .A(n22), .B(n3), .Z(\ab[9][16] ) );
  NR2 U92 ( .A(n22), .B(n4), .Z(\ab[9][15] ) );
  NR2 U93 ( .A(n22), .B(n5), .Z(\ab[9][14] ) );
  NR2 U94 ( .A(n22), .B(n6), .Z(\ab[9][13] ) );
  NR2 U95 ( .A(n22), .B(n7), .Z(\ab[9][12] ) );
  NR2 U96 ( .A(n22), .B(n8), .Z(\ab[9][11] ) );
  NR2 U97 ( .A(n22), .B(n9), .Z(\ab[9][10] ) );
  NR2 U98 ( .A(n22), .B(n19), .Z(\ab[9][0] ) );
  IV U99 ( .A(A[9]), .Z(n22) );
  NR2 U100 ( .A(n10), .B(n23), .Z(\ab[8][9] ) );
  NR2 U101 ( .A(n11), .B(n23), .Z(\ab[8][8] ) );
  NR2 U102 ( .A(n12), .B(n23), .Z(\ab[8][7] ) );
  NR2 U103 ( .A(n13), .B(n23), .Z(\ab[8][6] ) );
  NR2 U104 ( .A(n14), .B(n23), .Z(\ab[8][5] ) );
  NR2 U105 ( .A(n15), .B(n23), .Z(\ab[8][4] ) );
  NR2 U106 ( .A(n16), .B(n23), .Z(\ab[8][3] ) );
  NR2 U107 ( .A(n17), .B(n23), .Z(\ab[8][2] ) );
  NR2 U108 ( .A(n18), .B(n23), .Z(\ab[8][1] ) );
  NR2 U109 ( .A(n3), .B(n23), .Z(\ab[8][16] ) );
  NR2 U110 ( .A(n4), .B(n23), .Z(\ab[8][15] ) );
  NR2 U111 ( .A(n5), .B(n23), .Z(\ab[8][14] ) );
  NR2 U112 ( .A(n6), .B(n23), .Z(\ab[8][13] ) );
  NR2 U113 ( .A(n7), .B(n23), .Z(\ab[8][12] ) );
  NR2 U114 ( .A(n8), .B(n23), .Z(\ab[8][11] ) );
  NR2 U115 ( .A(n9), .B(n23), .Z(\ab[8][10] ) );
  NR2 U116 ( .A(n19), .B(n23), .Z(\ab[8][0] ) );
  IV U117 ( .A(A[8]), .Z(n23) );
  NR2 U118 ( .A(n10), .B(n24), .Z(\ab[7][9] ) );
  NR2 U119 ( .A(n11), .B(n24), .Z(\ab[7][8] ) );
  NR2 U120 ( .A(n12), .B(n24), .Z(\ab[7][7] ) );
  NR2 U121 ( .A(n13), .B(n24), .Z(\ab[7][6] ) );
  NR2 U122 ( .A(n14), .B(n24), .Z(\ab[7][5] ) );
  NR2 U123 ( .A(n15), .B(n24), .Z(\ab[7][4] ) );
  NR2 U124 ( .A(n16), .B(n24), .Z(\ab[7][3] ) );
  NR2 U125 ( .A(n17), .B(n24), .Z(\ab[7][2] ) );
  NR2 U126 ( .A(n18), .B(n24), .Z(\ab[7][1] ) );
  NR2 U127 ( .A(n3), .B(n24), .Z(\ab[7][16] ) );
  NR2 U128 ( .A(n4), .B(n24), .Z(\ab[7][15] ) );
  NR2 U129 ( .A(n5), .B(n24), .Z(\ab[7][14] ) );
  NR2 U130 ( .A(n6), .B(n24), .Z(\ab[7][13] ) );
  NR2 U131 ( .A(n7), .B(n24), .Z(\ab[7][12] ) );
  NR2 U132 ( .A(n8), .B(n24), .Z(\ab[7][11] ) );
  NR2 U133 ( .A(n9), .B(n24), .Z(\ab[7][10] ) );
  NR2 U134 ( .A(n19), .B(n24), .Z(\ab[7][0] ) );
  IV U135 ( .A(A[7]), .Z(n24) );
  NR2 U136 ( .A(n10), .B(n25), .Z(\ab[6][9] ) );
  NR2 U137 ( .A(n11), .B(n25), .Z(\ab[6][8] ) );
  NR2 U138 ( .A(n12), .B(n25), .Z(\ab[6][7] ) );
  NR2 U139 ( .A(n13), .B(n25), .Z(\ab[6][6] ) );
  NR2 U140 ( .A(n14), .B(n25), .Z(\ab[6][5] ) );
  NR2 U141 ( .A(n15), .B(n25), .Z(\ab[6][4] ) );
  NR2 U142 ( .A(n16), .B(n25), .Z(\ab[6][3] ) );
  NR2 U143 ( .A(n17), .B(n25), .Z(\ab[6][2] ) );
  NR2 U144 ( .A(n18), .B(n25), .Z(\ab[6][1] ) );
  NR2 U145 ( .A(n3), .B(n25), .Z(\ab[6][16] ) );
  NR2 U146 ( .A(n4), .B(n25), .Z(\ab[6][15] ) );
  NR2 U147 ( .A(n5), .B(n25), .Z(\ab[6][14] ) );
  NR2 U148 ( .A(n6), .B(n25), .Z(\ab[6][13] ) );
  NR2 U149 ( .A(n7), .B(n25), .Z(\ab[6][12] ) );
  NR2 U150 ( .A(n8), .B(n25), .Z(\ab[6][11] ) );
  NR2 U151 ( .A(n9), .B(n25), .Z(\ab[6][10] ) );
  NR2 U152 ( .A(n19), .B(n25), .Z(\ab[6][0] ) );
  IV U153 ( .A(A[6]), .Z(n25) );
  NR2 U154 ( .A(n10), .B(n26), .Z(\ab[5][9] ) );
  NR2 U155 ( .A(n11), .B(n26), .Z(\ab[5][8] ) );
  NR2 U156 ( .A(n12), .B(n26), .Z(\ab[5][7] ) );
  NR2 U157 ( .A(n13), .B(n26), .Z(\ab[5][6] ) );
  NR2 U158 ( .A(n14), .B(n26), .Z(\ab[5][5] ) );
  NR2 U159 ( .A(n15), .B(n26), .Z(\ab[5][4] ) );
  NR2 U160 ( .A(n16), .B(n26), .Z(\ab[5][3] ) );
  NR2 U161 ( .A(n17), .B(n26), .Z(\ab[5][2] ) );
  NR2 U162 ( .A(n18), .B(n26), .Z(\ab[5][1] ) );
  NR2 U163 ( .A(n3), .B(n26), .Z(\ab[5][16] ) );
  NR2 U164 ( .A(n4), .B(n26), .Z(\ab[5][15] ) );
  NR2 U165 ( .A(n5), .B(n26), .Z(\ab[5][14] ) );
  NR2 U166 ( .A(n6), .B(n26), .Z(\ab[5][13] ) );
  NR2 U167 ( .A(n7), .B(n26), .Z(\ab[5][12] ) );
  NR2 U168 ( .A(n8), .B(n26), .Z(\ab[5][11] ) );
  NR2 U169 ( .A(n9), .B(n26), .Z(\ab[5][10] ) );
  NR2 U170 ( .A(n19), .B(n26), .Z(\ab[5][0] ) );
  IV U171 ( .A(A[5]), .Z(n26) );
  NR2 U172 ( .A(n10), .B(n27), .Z(\ab[4][9] ) );
  NR2 U173 ( .A(n11), .B(n27), .Z(\ab[4][8] ) );
  NR2 U174 ( .A(n12), .B(n27), .Z(\ab[4][7] ) );
  NR2 U175 ( .A(n13), .B(n27), .Z(\ab[4][6] ) );
  NR2 U176 ( .A(n14), .B(n27), .Z(\ab[4][5] ) );
  NR2 U177 ( .A(n15), .B(n27), .Z(\ab[4][4] ) );
  NR2 U178 ( .A(n16), .B(n27), .Z(\ab[4][3] ) );
  NR2 U179 ( .A(n17), .B(n27), .Z(\ab[4][2] ) );
  NR2 U180 ( .A(n18), .B(n27), .Z(\ab[4][1] ) );
  NR2 U181 ( .A(n3), .B(n27), .Z(\ab[4][16] ) );
  NR2 U182 ( .A(n4), .B(n27), .Z(\ab[4][15] ) );
  NR2 U183 ( .A(n5), .B(n27), .Z(\ab[4][14] ) );
  NR2 U184 ( .A(n6), .B(n27), .Z(\ab[4][13] ) );
  NR2 U185 ( .A(n7), .B(n27), .Z(\ab[4][12] ) );
  NR2 U186 ( .A(n8), .B(n27), .Z(\ab[4][11] ) );
  NR2 U187 ( .A(n9), .B(n27), .Z(\ab[4][10] ) );
  NR2 U188 ( .A(n19), .B(n27), .Z(\ab[4][0] ) );
  IV U189 ( .A(A[4]), .Z(n27) );
  NR2 U190 ( .A(n10), .B(n28), .Z(\ab[3][9] ) );
  NR2 U191 ( .A(n11), .B(n28), .Z(\ab[3][8] ) );
  NR2 U192 ( .A(n12), .B(n28), .Z(\ab[3][7] ) );
  NR2 U193 ( .A(n13), .B(n28), .Z(\ab[3][6] ) );
  NR2 U194 ( .A(n14), .B(n28), .Z(\ab[3][5] ) );
  NR2 U195 ( .A(n15), .B(n28), .Z(\ab[3][4] ) );
  NR2 U196 ( .A(n16), .B(n28), .Z(\ab[3][3] ) );
  NR2 U197 ( .A(n17), .B(n28), .Z(\ab[3][2] ) );
  NR2 U198 ( .A(n18), .B(n28), .Z(\ab[3][1] ) );
  NR2 U199 ( .A(n3), .B(n28), .Z(\ab[3][16] ) );
  NR2 U200 ( .A(n4), .B(n28), .Z(\ab[3][15] ) );
  NR2 U201 ( .A(n5), .B(n28), .Z(\ab[3][14] ) );
  NR2 U202 ( .A(n6), .B(n28), .Z(\ab[3][13] ) );
  NR2 U203 ( .A(n7), .B(n28), .Z(\ab[3][12] ) );
  NR2 U204 ( .A(n8), .B(n28), .Z(\ab[3][11] ) );
  NR2 U205 ( .A(n9), .B(n28), .Z(\ab[3][10] ) );
  NR2 U206 ( .A(n19), .B(n28), .Z(\ab[3][0] ) );
  IV U207 ( .A(A[3]), .Z(n28) );
  NR2 U208 ( .A(n10), .B(n29), .Z(\ab[2][9] ) );
  NR2 U209 ( .A(n11), .B(n29), .Z(\ab[2][8] ) );
  NR2 U210 ( .A(n12), .B(n29), .Z(\ab[2][7] ) );
  NR2 U211 ( .A(n13), .B(n29), .Z(\ab[2][6] ) );
  NR2 U212 ( .A(n14), .B(n29), .Z(\ab[2][5] ) );
  NR2 U213 ( .A(n15), .B(n29), .Z(\ab[2][4] ) );
  NR2 U214 ( .A(n16), .B(n29), .Z(\ab[2][3] ) );
  NR2 U215 ( .A(n17), .B(n29), .Z(\ab[2][2] ) );
  NR2 U216 ( .A(n18), .B(n29), .Z(\ab[2][1] ) );
  NR2 U217 ( .A(n3), .B(n29), .Z(\ab[2][16] ) );
  NR2 U218 ( .A(n4), .B(n29), .Z(\ab[2][15] ) );
  NR2 U219 ( .A(n5), .B(n29), .Z(\ab[2][14] ) );
  NR2 U220 ( .A(n6), .B(n29), .Z(\ab[2][13] ) );
  NR2 U221 ( .A(n7), .B(n29), .Z(\ab[2][12] ) );
  NR2 U222 ( .A(n8), .B(n29), .Z(\ab[2][11] ) );
  NR2 U223 ( .A(n9), .B(n29), .Z(\ab[2][10] ) );
  NR2 U224 ( .A(n19), .B(n29), .Z(\ab[2][0] ) );
  IV U225 ( .A(A[2]), .Z(n29) );
  NR2 U226 ( .A(n10), .B(n30), .Z(\ab[1][9] ) );
  NR2 U227 ( .A(n11), .B(n30), .Z(\ab[1][8] ) );
  NR2 U228 ( .A(n12), .B(n30), .Z(\ab[1][7] ) );
  NR2 U229 ( .A(n13), .B(n30), .Z(\ab[1][6] ) );
  NR2 U230 ( .A(n14), .B(n30), .Z(\ab[1][5] ) );
  NR2 U231 ( .A(n15), .B(n30), .Z(\ab[1][4] ) );
  NR2 U232 ( .A(n16), .B(n30), .Z(\ab[1][3] ) );
  NR2 U233 ( .A(n17), .B(n30), .Z(\ab[1][2] ) );
  NR2 U234 ( .A(n3), .B(n30), .Z(\ab[1][16] ) );
  NR2 U235 ( .A(n4), .B(n30), .Z(\ab[1][15] ) );
  NR2 U236 ( .A(n5), .B(n30), .Z(\ab[1][14] ) );
  NR2 U237 ( .A(n6), .B(n30), .Z(\ab[1][13] ) );
  NR2 U238 ( .A(n7), .B(n30), .Z(\ab[1][12] ) );
  NR2 U239 ( .A(n8), .B(n30), .Z(\ab[1][11] ) );
  NR2 U240 ( .A(n9), .B(n30), .Z(\ab[1][10] ) );
  NR2 U241 ( .A(n10), .B(n31), .Z(\ab[14][9] ) );
  NR2 U242 ( .A(n11), .B(n31), .Z(\ab[14][8] ) );
  NR2 U243 ( .A(n12), .B(n31), .Z(\ab[14][7] ) );
  NR2 U244 ( .A(n13), .B(n31), .Z(\ab[14][6] ) );
  NR2 U245 ( .A(n14), .B(n31), .Z(\ab[14][5] ) );
  NR2 U246 ( .A(n15), .B(n31), .Z(\ab[14][4] ) );
  NR2 U247 ( .A(n16), .B(n31), .Z(\ab[14][3] ) );
  NR2 U248 ( .A(n17), .B(n31), .Z(\ab[14][2] ) );
  NR2 U249 ( .A(n18), .B(n31), .Z(\ab[14][1] ) );
  NR2 U250 ( .A(n3), .B(n31), .Z(\ab[14][16] ) );
  NR2 U251 ( .A(n4), .B(n31), .Z(\ab[14][15] ) );
  NR2 U252 ( .A(n5), .B(n31), .Z(\ab[14][14] ) );
  NR2 U253 ( .A(n6), .B(n31), .Z(\ab[14][13] ) );
  NR2 U254 ( .A(n7), .B(n31), .Z(\ab[14][12] ) );
  NR2 U255 ( .A(n8), .B(n31), .Z(\ab[14][11] ) );
  NR2 U256 ( .A(n9), .B(n31), .Z(\ab[14][10] ) );
  NR2 U257 ( .A(n19), .B(n31), .Z(\ab[14][0] ) );
  IV U258 ( .A(A[14]), .Z(n31) );
  NR2 U259 ( .A(n10), .B(n32), .Z(\ab[13][9] ) );
  NR2 U260 ( .A(n11), .B(n32), .Z(\ab[13][8] ) );
  NR2 U261 ( .A(n12), .B(n32), .Z(\ab[13][7] ) );
  NR2 U262 ( .A(n13), .B(n32), .Z(\ab[13][6] ) );
  NR2 U263 ( .A(n14), .B(n32), .Z(\ab[13][5] ) );
  NR2 U264 ( .A(n15), .B(n32), .Z(\ab[13][4] ) );
  NR2 U265 ( .A(n16), .B(n32), .Z(\ab[13][3] ) );
  NR2 U266 ( .A(n17), .B(n32), .Z(\ab[13][2] ) );
  NR2 U267 ( .A(n18), .B(n32), .Z(\ab[13][1] ) );
  NR2 U268 ( .A(n3), .B(n32), .Z(\ab[13][16] ) );
  NR2 U269 ( .A(n4), .B(n32), .Z(\ab[13][15] ) );
  NR2 U270 ( .A(n5), .B(n32), .Z(\ab[13][14] ) );
  NR2 U271 ( .A(n6), .B(n32), .Z(\ab[13][13] ) );
  NR2 U272 ( .A(n7), .B(n32), .Z(\ab[13][12] ) );
  NR2 U273 ( .A(n8), .B(n32), .Z(\ab[13][11] ) );
  NR2 U274 ( .A(n9), .B(n32), .Z(\ab[13][10] ) );
  NR2 U275 ( .A(n19), .B(n32), .Z(\ab[13][0] ) );
  IV U276 ( .A(A[13]), .Z(n32) );
  NR2 U277 ( .A(n10), .B(n33), .Z(\ab[12][9] ) );
  NR2 U278 ( .A(n11), .B(n33), .Z(\ab[12][8] ) );
  NR2 U279 ( .A(n12), .B(n33), .Z(\ab[12][7] ) );
  NR2 U280 ( .A(n13), .B(n33), .Z(\ab[12][6] ) );
  NR2 U281 ( .A(n14), .B(n33), .Z(\ab[12][5] ) );
  NR2 U282 ( .A(n15), .B(n33), .Z(\ab[12][4] ) );
  NR2 U283 ( .A(n16), .B(n33), .Z(\ab[12][3] ) );
  NR2 U284 ( .A(n17), .B(n33), .Z(\ab[12][2] ) );
  NR2 U285 ( .A(n18), .B(n33), .Z(\ab[12][1] ) );
  NR2 U286 ( .A(n3), .B(n33), .Z(\ab[12][16] ) );
  NR2 U287 ( .A(n4), .B(n33), .Z(\ab[12][15] ) );
  NR2 U288 ( .A(n5), .B(n33), .Z(\ab[12][14] ) );
  NR2 U289 ( .A(n6), .B(n33), .Z(\ab[12][13] ) );
  NR2 U290 ( .A(n7), .B(n33), .Z(\ab[12][12] ) );
  NR2 U291 ( .A(n8), .B(n33), .Z(\ab[12][11] ) );
  NR2 U292 ( .A(n9), .B(n33), .Z(\ab[12][10] ) );
  NR2 U293 ( .A(n19), .B(n33), .Z(\ab[12][0] ) );
  IV U294 ( .A(A[12]), .Z(n33) );
  NR2 U295 ( .A(n10), .B(n34), .Z(\ab[11][9] ) );
  NR2 U296 ( .A(n11), .B(n34), .Z(\ab[11][8] ) );
  NR2 U297 ( .A(n12), .B(n34), .Z(\ab[11][7] ) );
  NR2 U298 ( .A(n13), .B(n34), .Z(\ab[11][6] ) );
  NR2 U299 ( .A(n14), .B(n34), .Z(\ab[11][5] ) );
  NR2 U300 ( .A(n15), .B(n34), .Z(\ab[11][4] ) );
  NR2 U301 ( .A(n16), .B(n34), .Z(\ab[11][3] ) );
  NR2 U302 ( .A(n17), .B(n34), .Z(\ab[11][2] ) );
  NR2 U303 ( .A(n18), .B(n34), .Z(\ab[11][1] ) );
  NR2 U304 ( .A(n3), .B(n34), .Z(\ab[11][16] ) );
  NR2 U305 ( .A(n4), .B(n34), .Z(\ab[11][15] ) );
  NR2 U306 ( .A(n5), .B(n34), .Z(\ab[11][14] ) );
  NR2 U307 ( .A(n6), .B(n34), .Z(\ab[11][13] ) );
  NR2 U308 ( .A(n7), .B(n34), .Z(\ab[11][12] ) );
  NR2 U309 ( .A(n8), .B(n34), .Z(\ab[11][11] ) );
  NR2 U310 ( .A(n9), .B(n34), .Z(\ab[11][10] ) );
  NR2 U311 ( .A(n19), .B(n34), .Z(\ab[11][0] ) );
  IV U312 ( .A(A[11]), .Z(n34) );
  NR2 U313 ( .A(n10), .B(n35), .Z(\ab[10][9] ) );
  NR2 U314 ( .A(n11), .B(n35), .Z(\ab[10][8] ) );
  NR2 U315 ( .A(n12), .B(n35), .Z(\ab[10][7] ) );
  NR2 U316 ( .A(n13), .B(n35), .Z(\ab[10][6] ) );
  NR2 U317 ( .A(n14), .B(n35), .Z(\ab[10][5] ) );
  NR2 U318 ( .A(n15), .B(n35), .Z(\ab[10][4] ) );
  NR2 U319 ( .A(n16), .B(n35), .Z(\ab[10][3] ) );
  NR2 U320 ( .A(n17), .B(n35), .Z(\ab[10][2] ) );
  NR2 U321 ( .A(n18), .B(n35), .Z(\ab[10][1] ) );
  NR2 U322 ( .A(n3), .B(n35), .Z(\ab[10][16] ) );
  NR2 U323 ( .A(n4), .B(n35), .Z(\ab[10][15] ) );
  NR2 U324 ( .A(n5), .B(n35), .Z(\ab[10][14] ) );
  NR2 U325 ( .A(n6), .B(n35), .Z(\ab[10][13] ) );
  NR2 U326 ( .A(n7), .B(n35), .Z(\ab[10][12] ) );
  NR2 U327 ( .A(n8), .B(n35), .Z(\ab[10][11] ) );
  NR2 U328 ( .A(n9), .B(n35), .Z(\ab[10][10] ) );
  NR2 U329 ( .A(n19), .B(n35), .Z(\ab[10][0] ) );
  IV U330 ( .A(A[10]), .Z(n35) );
  NR2 U331 ( .A(n10), .B(n36), .Z(\ab[0][9] ) );
  NR2 U332 ( .A(n11), .B(n36), .Z(\ab[0][8] ) );
  NR2 U333 ( .A(n12), .B(n36), .Z(\ab[0][7] ) );
  NR2 U334 ( .A(n13), .B(n36), .Z(\ab[0][6] ) );
  NR2 U335 ( .A(n14), .B(n36), .Z(\ab[0][5] ) );
  NR2 U336 ( .A(n15), .B(n36), .Z(\ab[0][4] ) );
  NR2 U337 ( .A(n16), .B(n36), .Z(\ab[0][3] ) );
  NR2 U338 ( .A(n17), .B(n36), .Z(\ab[0][2] ) );
  NR2 U339 ( .A(n3), .B(n36), .Z(\ab[0][16] ) );
  NR2 U340 ( .A(n4), .B(n36), .Z(\ab[0][15] ) );
  NR2 U341 ( .A(n5), .B(n36), .Z(\ab[0][14] ) );
  NR2 U342 ( .A(n6), .B(n36), .Z(\ab[0][13] ) );
  NR2 U343 ( .A(n7), .B(n36), .Z(\ab[0][12] ) );
  NR2 U344 ( .A(n8), .B(n36), .Z(\ab[0][11] ) );
  NR2 U345 ( .A(n9), .B(n36), .Z(\ab[0][10] ) );
  IV U346 ( .A(A[0]), .Z(n36) );
  AN3 U347 ( .A(\ab[1][1] ), .B(B[0]), .C(A[0]), .Z(\CARRYB[1][0] ) );
  NR2 U348 ( .A(n30), .B(n18), .Z(\ab[1][1] ) );
  IV U349 ( .A(A[1]), .Z(n30) );
endmodule


module top_module ( clock, reset, X0_output, X1_output, valid );
  output [15:0] X0_output;
  output [15:0] X1_output;
  input clock, reset;
  output valid;
  wire   valid0, valid1, valid2, valid3, valid4, valid5, valid6, valid7,
         valid8, valid9, valid10, valid11, valid12, valid13, valid14, valid15,
         N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         N34, N50, N66, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365;
  wire   [31:0] taus_out_1;
  wire   [31:0] taus_out_0;
  wire   [47:0] LogIn;
  wire   [16:0] stage0;
  wire   [16:0] sqrt_out;
  wire   [16:0] stage1;
  wire   [16:0] stage2;
  wire   [16:0] stage3;
  wire   [16:0] stage4;
  wire   [16:0] stage5;
  wire   [16:0] stage6;
  wire   [16:0] sqrtOut;
  wire   [15:0] X0;
  wire   [15:0] X1;
  wire   [31:17] X0_reg;
  wire   [31:17] X1_reg;
  wire   [15:0] X01;
  wire   [15:0] X11;
  wire   [30:0] logarith_out;
  tri   clock;
  tri   [15:0] Angle;
  tri   [15:0] sin_out;
  tri   [15:0] cos_out;
  tri   n349;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;

  tausworthe_0 taus_gen ( .clock(clock), .re_set(reset), .tausout(taus_out_0)
         );
  tausworthe_1 taus_gen1 ( .clock(clock), .re_set(reset), .tausout(taus_out_1)
         );
  CORDIC codic_sin_cos ( .p1(clock), .p2(Angle), .p4({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p5(cos_out), .p6(sin_out) );
  Poly_Logarithm login ( .clock(clock), .reset(reset), .input_log(LogIn), 
        .output_log({logarith_out[30:1], SYNOPSYS_UNCONNECTED__0}) );
  Poly_sqrt sqrt1 ( .clock(clock), .reset(reset), .Datain({logarith_out[30:1], 
        1'b0}), .DataOut(sqrt_out) );
  top_module_DW02_mult_0 mult_79 ( .A(cos_out[14:0]), .B(sqrtOut), .TC(1'b0), 
        .PRODUCT({N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, 
        N22, N21, N20, SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17}) );
  top_module_DW02_mult_1 mult_78 ( .A(sin_out[14:0]), .B(sqrtOut), .TC(1'b0), 
        .PRODUCT({N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, 
        N6, N5, SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34}) );
  FD1 \Angle_reg[1]  ( .D(n364), .CP(clock), .Q(Angle[1]) );
  FD1 \Angle_reg[2]  ( .D(n363), .CP(clock), .Q(Angle[2]) );
  FD1 \Angle_reg[3]  ( .D(n350), .CP(clock), .Q(Angle[3]) );
  FD1 \Angle_reg[4]  ( .D(n354), .CP(clock), .Q(Angle[4]) );
  FD1 \Angle_reg[5]  ( .D(n357), .CP(clock), .Q(Angle[5]) );
  FD1 \Angle_reg[6]  ( .D(n360), .CP(clock), .Q(Angle[6]) );
  FD1 \Angle_reg[7]  ( .D(n351), .CP(clock), .Q(Angle[7]) );
  FD1 \Angle_reg[8]  ( .D(n355), .CP(clock), .Q(Angle[8]) );
  FD1 \Angle_reg[9]  ( .D(n358), .CP(clock), .Q(Angle[9]) );
  FD1 \Angle_reg[10]  ( .D(n361), .CP(clock), .Q(Angle[10]) );
  FD1 \Angle_reg[11]  ( .D(n352), .CP(clock), .Q(Angle[11]) );
  FD1 \Angle_reg[12]  ( .D(n356), .CP(clock), .Q(Angle[12]) );
  FD1 \Angle_reg[13]  ( .D(n359), .CP(clock), .Q(Angle[13]) );
  FD1 \Angle_reg[14]  ( .D(n362), .CP(clock), .Q(Angle[14]) );
  FD1 \Angle_reg[15]  ( .D(n353), .CP(clock), .Q(Angle[15]) );
  FDS2L \sqrtOut_reg[16]  ( .CR(1'b1), .D(stage6[16]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[16]) );
  FDS2L \sqrtOut_reg[15]  ( .CR(1'b1), .D(stage6[15]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[15]) );
  FDS2L \sqrtOut_reg[14]  ( .CR(1'b1), .D(stage6[14]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[14]) );
  FDS2L \sqrtOut_reg[13]  ( .CR(1'b1), .D(stage6[13]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[13]) );
  FDS2L \sqrtOut_reg[12]  ( .CR(1'b1), .D(stage6[12]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[12]) );
  FDS2L \sqrtOut_reg[11]  ( .CR(1'b1), .D(stage6[11]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[11]) );
  FDS2L \sqrtOut_reg[10]  ( .CR(1'b1), .D(stage6[10]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[10]) );
  FDS2L \sqrtOut_reg[9]  ( .CR(1'b1), .D(stage6[9]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[9]) );
  FDS2L \sqrtOut_reg[8]  ( .CR(1'b1), .D(stage6[8]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[8]) );
  FDS2L \sqrtOut_reg[7]  ( .CR(1'b1), .D(stage6[7]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[7]) );
  FDS2L \sqrtOut_reg[6]  ( .CR(1'b1), .D(stage6[6]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[6]) );
  FDS2L \sqrtOut_reg[5]  ( .CR(1'b1), .D(stage6[5]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[5]) );
  FDS2L \sqrtOut_reg[4]  ( .CR(1'b1), .D(stage6[4]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[4]) );
  FDS2L \sqrtOut_reg[3]  ( .CR(1'b1), .D(stage6[3]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[3]) );
  FDS2L \sqrtOut_reg[2]  ( .CR(1'b1), .D(stage6[2]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[2]) );
  FDS2L \sqrtOut_reg[1]  ( .CR(1'b1), .D(stage6[1]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[1]) );
  FDS2L \sqrtOut_reg[0]  ( .CR(1'b1), .D(stage6[0]), .LD(n365), .CP(clock), 
        .Q(sqrtOut[0]) );
  FDS2L \Angle_reg[0]  ( .CR(1'b1), .D(taus_out_0[0]), .LD(n365), .CP(clock), 
        .Q(Angle[0]) );
  FDS2 valid_reg ( .CR(valid15), .D(n365), .CP(clock), .Q(valid) );
  FDS2L \X1_output_reg[15]  ( .CR(1'b1), .D(X11[15]), .LD(n365), .CP(clock), 
        .Q(X1_output[15]) );
  FDS2L \X1_output_reg[14]  ( .CR(1'b1), .D(X11[14]), .LD(n365), .CP(clock), 
        .Q(X1_output[14]) );
  FDS2L \X1_output_reg[13]  ( .CR(1'b1), .D(X11[13]), .LD(n365), .CP(clock), 
        .Q(X1_output[13]) );
  FDS2L \X1_output_reg[12]  ( .CR(1'b1), .D(X11[12]), .LD(n365), .CP(clock), 
        .Q(X1_output[12]) );
  FDS2L \X1_output_reg[11]  ( .CR(1'b1), .D(X11[11]), .LD(n365), .CP(clock), 
        .Q(X1_output[11]) );
  FDS2L \X1_output_reg[10]  ( .CR(1'b1), .D(X11[10]), .LD(n365), .CP(clock), 
        .Q(X1_output[10]) );
  FDS2L \X1_output_reg[9]  ( .CR(1'b1), .D(X11[9]), .LD(n365), .CP(clock), .Q(
        X1_output[9]) );
  FDS2L \X1_output_reg[8]  ( .CR(1'b1), .D(X11[8]), .LD(n365), .CP(clock), .Q(
        X1_output[8]) );
  FDS2L \X1_output_reg[7]  ( .CR(1'b1), .D(X11[7]), .LD(n365), .CP(clock), .Q(
        X1_output[7]) );
  FDS2L \X1_output_reg[6]  ( .CR(1'b1), .D(X11[6]), .LD(n365), .CP(clock), .Q(
        X1_output[6]) );
  FDS2L \X1_output_reg[5]  ( .CR(1'b1), .D(X11[5]), .LD(n365), .CP(clock), .Q(
        X1_output[5]) );
  FDS2L \X1_output_reg[4]  ( .CR(1'b1), .D(X11[4]), .LD(n365), .CP(clock), .Q(
        X1_output[4]) );
  FDS2L \X1_output_reg[3]  ( .CR(1'b1), .D(X11[3]), .LD(n365), .CP(clock), .Q(
        X1_output[3]) );
  FDS2L \X1_output_reg[2]  ( .CR(1'b1), .D(X11[2]), .LD(n365), .CP(clock), .Q(
        X1_output[2]) );
  FDS2L \X1_output_reg[1]  ( .CR(1'b1), .D(X11[1]), .LD(n365), .CP(clock), .Q(
        X1_output[1]) );
  FDS2L \X1_output_reg[0]  ( .CR(1'b1), .D(X11[0]), .LD(n365), .CP(clock), .Q(
        X1_output[0]) );
  FDS2L \X0_output_reg[15]  ( .CR(1'b1), .D(X01[15]), .LD(n365), .CP(clock), 
        .Q(X0_output[15]) );
  FDS2L \X0_output_reg[14]  ( .CR(1'b1), .D(X01[14]), .LD(n365), .CP(clock), 
        .Q(X0_output[14]) );
  FDS2L \X0_output_reg[13]  ( .CR(1'b1), .D(X01[13]), .LD(n365), .CP(clock), 
        .Q(X0_output[13]) );
  FDS2L \X0_output_reg[12]  ( .CR(1'b1), .D(X01[12]), .LD(n365), .CP(clock), 
        .Q(X0_output[12]) );
  FDS2L \X0_output_reg[11]  ( .CR(1'b1), .D(X01[11]), .LD(n365), .CP(clock), 
        .Q(X0_output[11]) );
  FDS2L \X0_output_reg[10]  ( .CR(1'b1), .D(X01[10]), .LD(n365), .CP(clock), 
        .Q(X0_output[10]) );
  FDS2L \X0_output_reg[9]  ( .CR(1'b1), .D(X01[9]), .LD(n365), .CP(clock), .Q(
        X0_output[9]) );
  FDS2L \X0_output_reg[8]  ( .CR(1'b1), .D(X01[8]), .LD(n365), .CP(clock), .Q(
        X0_output[8]) );
  FDS2L \X0_output_reg[7]  ( .CR(1'b1), .D(X01[7]), .LD(n365), .CP(clock), .Q(
        X0_output[7]) );
  FDS2L \X0_output_reg[6]  ( .CR(1'b1), .D(X01[6]), .LD(n365), .CP(clock), .Q(
        X0_output[6]) );
  FDS2L \X0_output_reg[5]  ( .CR(1'b1), .D(X01[5]), .LD(n365), .CP(clock), .Q(
        X0_output[5]) );
  FDS2L \X0_output_reg[4]  ( .CR(1'b1), .D(X01[4]), .LD(n365), .CP(clock), .Q(
        X0_output[4]) );
  FDS2L \X0_output_reg[3]  ( .CR(1'b1), .D(X01[3]), .LD(n365), .CP(clock), .Q(
        X0_output[3]) );
  FDS2L \X0_output_reg[2]  ( .CR(1'b1), .D(X01[2]), .LD(n365), .CP(clock), .Q(
        X0_output[2]) );
  FDS2L \X0_output_reg[1]  ( .CR(1'b1), .D(X01[1]), .LD(n365), .CP(clock), .Q(
        X0_output[1]) );
  FDS2L \X0_output_reg[0]  ( .CR(1'b1), .D(X01[0]), .LD(n365), .CP(clock), .Q(
        X0_output[0]) );
  FD1 valid0_reg ( .D(n365), .CP(clock), .Q(valid0) );
  FDS2 valid1_reg ( .CR(valid0), .D(n365), .CP(clock), .Q(valid1) );
  FDS2 valid2_reg ( .CR(valid1), .D(n365), .CP(clock), .Q(valid2) );
  FDS2 valid3_reg ( .CR(valid2), .D(n365), .CP(clock), .Q(valid3) );
  FDS2 valid4_reg ( .CR(valid3), .D(n365), .CP(clock), .Q(valid4) );
  FDS2 valid5_reg ( .CR(valid4), .D(n365), .CP(clock), .Q(valid5) );
  FDS2 valid6_reg ( .CR(valid5), .D(n365), .CP(clock), .Q(valid6) );
  FDS2 valid7_reg ( .CR(valid6), .D(n365), .CP(clock), .Q(valid7) );
  FDS2 valid8_reg ( .CR(valid7), .D(n365), .CP(clock), .Q(valid8) );
  FDS2 valid9_reg ( .CR(valid8), .D(n365), .CP(clock), .Q(valid9) );
  FDS2 valid10_reg ( .CR(valid9), .D(n365), .CP(clock), .Q(valid10) );
  FDS2 valid11_reg ( .CR(valid10), .D(n365), .CP(clock), .Q(valid11) );
  FDS2 valid12_reg ( .CR(valid11), .D(n365), .CP(clock), .Q(valid12) );
  FDS2 valid13_reg ( .CR(valid12), .D(n365), .CP(clock), .Q(valid13) );
  FDS2 valid14_reg ( .CR(valid13), .D(n365), .CP(clock), .Q(valid14) );
  FDS2 valid15_reg ( .CR(valid14), .D(n365), .CP(clock), .Q(valid15) );
  FDS2L \LogIn_reg[16]  ( .CR(1'b1), .D(taus_out_1[0]), .LD(n365), .CP(clock), 
        .Q(LogIn[16]) );
  FDS2L \LogIn_reg[17]  ( .CR(1'b1), .D(taus_out_1[1]), .LD(n365), .CP(clock), 
        .Q(LogIn[17]) );
  FDS2L \LogIn_reg[18]  ( .CR(1'b1), .D(taus_out_1[2]), .LD(n365), .CP(clock), 
        .Q(LogIn[18]) );
  FDS2L \LogIn_reg[19]  ( .CR(1'b1), .D(taus_out_1[3]), .LD(n365), .CP(clock), 
        .Q(LogIn[19]) );
  FDS2L \LogIn_reg[20]  ( .CR(1'b1), .D(taus_out_1[4]), .LD(n365), .CP(clock), 
        .Q(LogIn[20]) );
  FDS2L \LogIn_reg[21]  ( .CR(1'b1), .D(taus_out_1[5]), .LD(n365), .CP(clock), 
        .Q(LogIn[21]) );
  FDS2L \LogIn_reg[22]  ( .CR(1'b1), .D(taus_out_1[6]), .LD(n365), .CP(clock), 
        .Q(LogIn[22]) );
  FDS2L \LogIn_reg[23]  ( .CR(1'b1), .D(taus_out_1[7]), .LD(n365), .CP(clock), 
        .Q(LogIn[23]) );
  FDS2L \LogIn_reg[24]  ( .CR(1'b1), .D(taus_out_1[8]), .LD(n365), .CP(clock), 
        .Q(LogIn[24]) );
  FDS2L \LogIn_reg[25]  ( .CR(1'b1), .D(taus_out_1[9]), .LD(n365), .CP(clock), 
        .Q(LogIn[25]) );
  FDS2L \LogIn_reg[26]  ( .CR(1'b1), .D(taus_out_1[10]), .LD(n365), .CP(clock), 
        .Q(LogIn[26]) );
  FDS2L \LogIn_reg[27]  ( .CR(1'b1), .D(taus_out_1[11]), .LD(n365), .CP(clock), 
        .Q(LogIn[27]) );
  FDS2L \LogIn_reg[28]  ( .CR(1'b1), .D(taus_out_1[12]), .LD(n365), .CP(clock), 
        .Q(LogIn[28]) );
  FDS2L \LogIn_reg[29]  ( .CR(1'b1), .D(taus_out_1[13]), .LD(n365), .CP(clock), 
        .Q(LogIn[29]) );
  FDS2L \LogIn_reg[30]  ( .CR(1'b1), .D(taus_out_1[14]), .LD(n365), .CP(clock), 
        .Q(LogIn[30]) );
  FDS2L \LogIn_reg[31]  ( .CR(1'b1), .D(taus_out_1[15]), .LD(n365), .CP(clock), 
        .Q(LogIn[31]) );
  FDS2L \LogIn_reg[32]  ( .CR(1'b1), .D(taus_out_1[16]), .LD(n365), .CP(clock), 
        .Q(LogIn[32]) );
  FDS2L \LogIn_reg[33]  ( .CR(1'b1), .D(taus_out_1[17]), .LD(n365), .CP(clock), 
        .Q(LogIn[33]) );
  FDS2L \LogIn_reg[34]  ( .CR(1'b1), .D(taus_out_1[18]), .LD(n365), .CP(clock), 
        .Q(LogIn[34]) );
  FDS2L \LogIn_reg[35]  ( .CR(1'b1), .D(taus_out_1[19]), .LD(n365), .CP(clock), 
        .Q(LogIn[35]) );
  FDS2L \LogIn_reg[36]  ( .CR(1'b1), .D(taus_out_1[20]), .LD(n365), .CP(clock), 
        .Q(LogIn[36]) );
  FDS2L \LogIn_reg[37]  ( .CR(1'b1), .D(taus_out_1[21]), .LD(n365), .CP(clock), 
        .Q(LogIn[37]) );
  FDS2L \LogIn_reg[38]  ( .CR(1'b1), .D(taus_out_1[22]), .LD(n365), .CP(clock), 
        .Q(LogIn[38]) );
  FDS2L \LogIn_reg[39]  ( .CR(1'b1), .D(taus_out_1[23]), .LD(n365), .CP(clock), 
        .Q(LogIn[39]) );
  FDS2L \LogIn_reg[40]  ( .CR(1'b1), .D(taus_out_1[24]), .LD(n365), .CP(clock), 
        .Q(LogIn[40]) );
  FDS2L \LogIn_reg[41]  ( .CR(1'b1), .D(taus_out_1[25]), .LD(n365), .CP(clock), 
        .Q(LogIn[41]) );
  FDS2L \LogIn_reg[42]  ( .CR(1'b1), .D(taus_out_1[26]), .LD(n365), .CP(clock), 
        .Q(LogIn[42]) );
  FDS2L \LogIn_reg[43]  ( .CR(1'b1), .D(taus_out_1[27]), .LD(n365), .CP(clock), 
        .Q(LogIn[43]) );
  FDS2L \LogIn_reg[44]  ( .CR(1'b1), .D(taus_out_1[28]), .LD(n365), .CP(clock), 
        .Q(LogIn[44]) );
  FDS2L \LogIn_reg[45]  ( .CR(1'b1), .D(taus_out_1[29]), .LD(n365), .CP(clock), 
        .Q(LogIn[45]) );
  FDS2L \LogIn_reg[46]  ( .CR(1'b1), .D(taus_out_1[30]), .LD(n365), .CP(clock), 
        .Q(LogIn[46]) );
  FDS2L \LogIn_reg[47]  ( .CR(1'b1), .D(taus_out_1[31]), .LD(n365), .CP(clock), 
        .Q(LogIn[47]) );
  FDS2L \LogIn_reg[0]  ( .CR(1'b1), .D(taus_out_0[16]), .LD(n365), .CP(clock), 
        .Q(LogIn[0]) );
  FDS2L \LogIn_reg[1]  ( .CR(1'b1), .D(taus_out_0[17]), .LD(n365), .CP(clock), 
        .Q(LogIn[1]) );
  FDS2L \LogIn_reg[2]  ( .CR(1'b1), .D(taus_out_0[18]), .LD(n365), .CP(clock), 
        .Q(LogIn[2]) );
  FDS2L \LogIn_reg[3]  ( .CR(1'b1), .D(taus_out_0[19]), .LD(n365), .CP(clock), 
        .Q(LogIn[3]) );
  FDS2L \LogIn_reg[4]  ( .CR(1'b1), .D(taus_out_0[20]), .LD(n365), .CP(clock), 
        .Q(LogIn[4]) );
  FDS2L \LogIn_reg[5]  ( .CR(1'b1), .D(taus_out_0[21]), .LD(n365), .CP(clock), 
        .Q(LogIn[5]) );
  FDS2L \LogIn_reg[6]  ( .CR(1'b1), .D(taus_out_0[22]), .LD(n365), .CP(clock), 
        .Q(LogIn[6]) );
  FDS2L \LogIn_reg[7]  ( .CR(1'b1), .D(taus_out_0[23]), .LD(n365), .CP(clock), 
        .Q(LogIn[7]) );
  FDS2L \LogIn_reg[8]  ( .CR(1'b1), .D(taus_out_0[24]), .LD(n365), .CP(clock), 
        .Q(LogIn[8]) );
  FDS2L \LogIn_reg[9]  ( .CR(1'b1), .D(taus_out_0[25]), .LD(n365), .CP(clock), 
        .Q(LogIn[9]) );
  FDS2L \LogIn_reg[10]  ( .CR(1'b1), .D(taus_out_0[26]), .LD(n365), .CP(clock), 
        .Q(LogIn[10]) );
  FDS2L \LogIn_reg[11]  ( .CR(1'b1), .D(taus_out_0[27]), .LD(n365), .CP(clock), 
        .Q(LogIn[11]) );
  FDS2L \LogIn_reg[12]  ( .CR(1'b1), .D(taus_out_0[28]), .LD(n365), .CP(clock), 
        .Q(LogIn[12]) );
  FDS2L \LogIn_reg[13]  ( .CR(1'b1), .D(taus_out_0[29]), .LD(n365), .CP(clock), 
        .Q(LogIn[13]) );
  FDS2L \LogIn_reg[14]  ( .CR(1'b1), .D(taus_out_0[30]), .LD(n365), .CP(clock), 
        .Q(LogIn[14]) );
  FDS2L \LogIn_reg[15]  ( .CR(1'b1), .D(taus_out_0[31]), .LD(n365), .CP(clock), 
        .Q(LogIn[15]) );
  FDS2L \stage0_reg[16]  ( .CR(1'b1), .D(sqrt_out[16]), .LD(n365), .CP(clock), 
        .Q(stage0[16]) );
  FDS2L \stage0_reg[15]  ( .CR(1'b1), .D(sqrt_out[15]), .LD(n365), .CP(clock), 
        .Q(stage0[15]) );
  FDS2L \stage0_reg[14]  ( .CR(1'b1), .D(sqrt_out[14]), .LD(n365), .CP(clock), 
        .Q(stage0[14]) );
  FDS2L \stage0_reg[13]  ( .CR(1'b1), .D(sqrt_out[13]), .LD(n365), .CP(clock), 
        .Q(stage0[13]) );
  FDS2L \stage0_reg[12]  ( .CR(1'b1), .D(sqrt_out[12]), .LD(n365), .CP(clock), 
        .Q(stage0[12]) );
  FDS2L \stage0_reg[11]  ( .CR(1'b1), .D(sqrt_out[11]), .LD(n365), .CP(clock), 
        .Q(stage0[11]) );
  FDS2L \stage0_reg[10]  ( .CR(1'b1), .D(sqrt_out[10]), .LD(n365), .CP(clock), 
        .Q(stage0[10]) );
  FDS2L \stage0_reg[9]  ( .CR(1'b1), .D(sqrt_out[9]), .LD(n365), .CP(clock), 
        .Q(stage0[9]) );
  FDS2L \stage0_reg[8]  ( .CR(1'b1), .D(sqrt_out[8]), .LD(n365), .CP(clock), 
        .Q(stage0[8]) );
  FDS2L \stage0_reg[7]  ( .CR(1'b1), .D(sqrt_out[7]), .LD(n365), .CP(clock), 
        .Q(stage0[7]) );
  FDS2L \stage0_reg[6]  ( .CR(1'b1), .D(sqrt_out[6]), .LD(n365), .CP(clock), 
        .Q(stage0[6]) );
  FDS2L \stage0_reg[5]  ( .CR(1'b1), .D(sqrt_out[5]), .LD(n365), .CP(clock), 
        .Q(stage0[5]) );
  FDS2L \stage0_reg[4]  ( .CR(1'b1), .D(sqrt_out[4]), .LD(n365), .CP(clock), 
        .Q(stage0[4]) );
  FDS2L \stage0_reg[3]  ( .CR(1'b1), .D(sqrt_out[3]), .LD(n365), .CP(clock), 
        .Q(stage0[3]) );
  FDS2L \stage0_reg[2]  ( .CR(1'b1), .D(sqrt_out[2]), .LD(n365), .CP(clock), 
        .Q(stage0[2]) );
  FDS2L \stage0_reg[1]  ( .CR(1'b1), .D(sqrt_out[1]), .LD(n365), .CP(clock), 
        .Q(stage0[1]) );
  FDS2L \stage0_reg[0]  ( .CR(1'b1), .D(sqrt_out[0]), .LD(n365), .CP(clock), 
        .Q(stage0[0]) );
  FDS2L \stage1_reg[16]  ( .CR(1'b1), .D(stage0[16]), .LD(n365), .CP(clock), 
        .Q(stage1[16]) );
  FDS2L \stage1_reg[15]  ( .CR(1'b1), .D(stage0[15]), .LD(n365), .CP(clock), 
        .Q(stage1[15]) );
  FDS2L \stage1_reg[14]  ( .CR(1'b1), .D(stage0[14]), .LD(n365), .CP(clock), 
        .Q(stage1[14]) );
  FDS2L \stage1_reg[13]  ( .CR(1'b1), .D(stage0[13]), .LD(n365), .CP(clock), 
        .Q(stage1[13]) );
  FDS2L \stage1_reg[12]  ( .CR(1'b1), .D(stage0[12]), .LD(n365), .CP(clock), 
        .Q(stage1[12]) );
  FDS2L \stage1_reg[11]  ( .CR(1'b1), .D(stage0[11]), .LD(n365), .CP(clock), 
        .Q(stage1[11]) );
  FDS2L \stage1_reg[10]  ( .CR(1'b1), .D(stage0[10]), .LD(n365), .CP(clock), 
        .Q(stage1[10]) );
  FDS2L \stage1_reg[9]  ( .CR(1'b1), .D(stage0[9]), .LD(n365), .CP(clock), .Q(
        stage1[9]) );
  FDS2L \stage1_reg[8]  ( .CR(1'b1), .D(stage0[8]), .LD(n365), .CP(clock), .Q(
        stage1[8]) );
  FDS2L \stage1_reg[7]  ( .CR(1'b1), .D(stage0[7]), .LD(n365), .CP(clock), .Q(
        stage1[7]) );
  FDS2L \stage1_reg[6]  ( .CR(1'b1), .D(stage0[6]), .LD(n365), .CP(clock), .Q(
        stage1[6]) );
  FDS2L \stage1_reg[5]  ( .CR(1'b1), .D(stage0[5]), .LD(n365), .CP(clock), .Q(
        stage1[5]) );
  FDS2L \stage1_reg[4]  ( .CR(1'b1), .D(stage0[4]), .LD(n365), .CP(clock), .Q(
        stage1[4]) );
  FDS2L \stage1_reg[3]  ( .CR(1'b1), .D(stage0[3]), .LD(n365), .CP(clock), .Q(
        stage1[3]) );
  FDS2L \stage1_reg[2]  ( .CR(1'b1), .D(stage0[2]), .LD(n365), .CP(clock), .Q(
        stage1[2]) );
  FDS2L \stage1_reg[1]  ( .CR(1'b1), .D(stage0[1]), .LD(n365), .CP(clock), .Q(
        stage1[1]) );
  FDS2L \stage1_reg[0]  ( .CR(1'b1), .D(stage0[0]), .LD(n365), .CP(clock), .Q(
        stage1[0]) );
  FDS2L \stage2_reg[16]  ( .CR(1'b1), .D(stage1[16]), .LD(n365), .CP(clock), 
        .Q(stage2[16]) );
  FDS2L \stage2_reg[15]  ( .CR(1'b1), .D(stage1[15]), .LD(n365), .CP(clock), 
        .Q(stage2[15]) );
  FDS2L \stage2_reg[14]  ( .CR(1'b1), .D(stage1[14]), .LD(n365), .CP(clock), 
        .Q(stage2[14]) );
  FDS2L \stage2_reg[13]  ( .CR(1'b1), .D(stage1[13]), .LD(n365), .CP(clock), 
        .Q(stage2[13]) );
  FDS2L \stage2_reg[12]  ( .CR(1'b1), .D(stage1[12]), .LD(n365), .CP(clock), 
        .Q(stage2[12]) );
  FDS2L \stage2_reg[11]  ( .CR(1'b1), .D(stage1[11]), .LD(n365), .CP(clock), 
        .Q(stage2[11]) );
  FDS2L \stage2_reg[10]  ( .CR(1'b1), .D(stage1[10]), .LD(n365), .CP(clock), 
        .Q(stage2[10]) );
  FDS2L \stage2_reg[9]  ( .CR(1'b1), .D(stage1[9]), .LD(n365), .CP(clock), .Q(
        stage2[9]) );
  FDS2L \stage2_reg[8]  ( .CR(1'b1), .D(stage1[8]), .LD(n365), .CP(clock), .Q(
        stage2[8]) );
  FDS2L \stage2_reg[7]  ( .CR(1'b1), .D(stage1[7]), .LD(n365), .CP(clock), .Q(
        stage2[7]) );
  FDS2L \stage2_reg[6]  ( .CR(1'b1), .D(stage1[6]), .LD(n365), .CP(clock), .Q(
        stage2[6]) );
  FDS2L \stage2_reg[5]  ( .CR(1'b1), .D(stage1[5]), .LD(n365), .CP(clock), .Q(
        stage2[5]) );
  FDS2L \stage2_reg[4]  ( .CR(1'b1), .D(stage1[4]), .LD(n365), .CP(clock), .Q(
        stage2[4]) );
  FDS2L \stage2_reg[3]  ( .CR(1'b1), .D(stage1[3]), .LD(n365), .CP(clock), .Q(
        stage2[3]) );
  FDS2L \stage2_reg[2]  ( .CR(1'b1), .D(stage1[2]), .LD(n365), .CP(clock), .Q(
        stage2[2]) );
  FDS2L \stage2_reg[1]  ( .CR(1'b1), .D(stage1[1]), .LD(n365), .CP(clock), .Q(
        stage2[1]) );
  FDS2L \stage2_reg[0]  ( .CR(1'b1), .D(stage1[0]), .LD(n365), .CP(clock), .Q(
        stage2[0]) );
  FDS2L \stage3_reg[16]  ( .CR(1'b1), .D(stage2[16]), .LD(n365), .CP(clock), 
        .Q(stage3[16]) );
  FDS2L \stage3_reg[15]  ( .CR(1'b1), .D(stage2[15]), .LD(n365), .CP(clock), 
        .Q(stage3[15]) );
  FDS2L \stage3_reg[14]  ( .CR(1'b1), .D(stage2[14]), .LD(n365), .CP(clock), 
        .Q(stage3[14]) );
  FDS2L \stage3_reg[13]  ( .CR(1'b1), .D(stage2[13]), .LD(n365), .CP(clock), 
        .Q(stage3[13]) );
  FDS2L \stage3_reg[12]  ( .CR(1'b1), .D(stage2[12]), .LD(n365), .CP(clock), 
        .Q(stage3[12]) );
  FDS2L \stage3_reg[11]  ( .CR(1'b1), .D(stage2[11]), .LD(n365), .CP(clock), 
        .Q(stage3[11]) );
  FDS2L \stage3_reg[10]  ( .CR(1'b1), .D(stage2[10]), .LD(n365), .CP(clock), 
        .Q(stage3[10]) );
  FDS2L \stage3_reg[9]  ( .CR(1'b1), .D(stage2[9]), .LD(n365), .CP(clock), .Q(
        stage3[9]) );
  FDS2L \stage3_reg[8]  ( .CR(1'b1), .D(stage2[8]), .LD(n365), .CP(clock), .Q(
        stage3[8]) );
  FDS2L \stage3_reg[7]  ( .CR(1'b1), .D(stage2[7]), .LD(n365), .CP(clock), .Q(
        stage3[7]) );
  FDS2L \stage3_reg[6]  ( .CR(1'b1), .D(stage2[6]), .LD(n365), .CP(clock), .Q(
        stage3[6]) );
  FDS2L \stage3_reg[5]  ( .CR(1'b1), .D(stage2[5]), .LD(n365), .CP(clock), .Q(
        stage3[5]) );
  FDS2L \stage3_reg[4]  ( .CR(1'b1), .D(stage2[4]), .LD(n365), .CP(clock), .Q(
        stage3[4]) );
  FDS2L \stage3_reg[3]  ( .CR(1'b1), .D(stage2[3]), .LD(n365), .CP(clock), .Q(
        stage3[3]) );
  FDS2L \stage3_reg[2]  ( .CR(1'b1), .D(stage2[2]), .LD(n365), .CP(clock), .Q(
        stage3[2]) );
  FDS2L \stage3_reg[1]  ( .CR(1'b1), .D(stage2[1]), .LD(n365), .CP(clock), .Q(
        stage3[1]) );
  FDS2L \stage3_reg[0]  ( .CR(1'b1), .D(stage2[0]), .LD(n365), .CP(clock), .Q(
        stage3[0]) );
  FDS2L \stage4_reg[16]  ( .CR(1'b1), .D(stage3[16]), .LD(n365), .CP(clock), 
        .Q(stage4[16]) );
  FDS2L \stage4_reg[15]  ( .CR(1'b1), .D(stage3[15]), .LD(n365), .CP(clock), 
        .Q(stage4[15]) );
  FDS2L \stage4_reg[14]  ( .CR(1'b1), .D(stage3[14]), .LD(n365), .CP(clock), 
        .Q(stage4[14]) );
  FDS2L \stage4_reg[13]  ( .CR(1'b1), .D(stage3[13]), .LD(n365), .CP(clock), 
        .Q(stage4[13]) );
  FDS2L \stage4_reg[12]  ( .CR(1'b1), .D(stage3[12]), .LD(n365), .CP(clock), 
        .Q(stage4[12]) );
  FDS2L \stage4_reg[11]  ( .CR(1'b1), .D(stage3[11]), .LD(n365), .CP(clock), 
        .Q(stage4[11]) );
  FDS2L \stage4_reg[10]  ( .CR(1'b1), .D(stage3[10]), .LD(n365), .CP(clock), 
        .Q(stage4[10]) );
  FDS2L \stage4_reg[9]  ( .CR(1'b1), .D(stage3[9]), .LD(n365), .CP(clock), .Q(
        stage4[9]) );
  FDS2L \stage4_reg[8]  ( .CR(1'b1), .D(stage3[8]), .LD(n365), .CP(clock), .Q(
        stage4[8]) );
  FDS2L \stage4_reg[7]  ( .CR(1'b1), .D(stage3[7]), .LD(n365), .CP(clock), .Q(
        stage4[7]) );
  FDS2L \stage4_reg[6]  ( .CR(1'b1), .D(stage3[6]), .LD(n365), .CP(clock), .Q(
        stage4[6]) );
  FDS2L \stage4_reg[5]  ( .CR(1'b1), .D(stage3[5]), .LD(n365), .CP(clock), .Q(
        stage4[5]) );
  FDS2L \stage4_reg[4]  ( .CR(1'b1), .D(stage3[4]), .LD(n365), .CP(clock), .Q(
        stage4[4]) );
  FDS2L \stage4_reg[3]  ( .CR(1'b1), .D(stage3[3]), .LD(n365), .CP(clock), .Q(
        stage4[3]) );
  FDS2L \stage4_reg[2]  ( .CR(1'b1), .D(stage3[2]), .LD(n365), .CP(clock), .Q(
        stage4[2]) );
  FDS2L \stage4_reg[1]  ( .CR(1'b1), .D(stage3[1]), .LD(n365), .CP(clock), .Q(
        stage4[1]) );
  FDS2L \stage4_reg[0]  ( .CR(1'b1), .D(stage3[0]), .LD(n365), .CP(clock), .Q(
        stage4[0]) );
  FDS2L \stage5_reg[16]  ( .CR(1'b1), .D(stage4[16]), .LD(n365), .CP(clock), 
        .Q(stage5[16]) );
  FDS2L \stage5_reg[15]  ( .CR(1'b1), .D(stage4[15]), .LD(n365), .CP(clock), 
        .Q(stage5[15]) );
  FDS2L \stage5_reg[14]  ( .CR(1'b1), .D(stage4[14]), .LD(n365), .CP(clock), 
        .Q(stage5[14]) );
  FDS2L \stage5_reg[13]  ( .CR(1'b1), .D(stage4[13]), .LD(n365), .CP(clock), 
        .Q(stage5[13]) );
  FDS2L \stage5_reg[12]  ( .CR(1'b1), .D(stage4[12]), .LD(n365), .CP(clock), 
        .Q(stage5[12]) );
  FDS2L \stage5_reg[11]  ( .CR(1'b1), .D(stage4[11]), .LD(n365), .CP(clock), 
        .Q(stage5[11]) );
  FDS2L \stage5_reg[10]  ( .CR(1'b1), .D(stage4[10]), .LD(n365), .CP(clock), 
        .Q(stage5[10]) );
  FDS2L \stage5_reg[9]  ( .CR(1'b1), .D(stage4[9]), .LD(n365), .CP(clock), .Q(
        stage5[9]) );
  FDS2L \stage5_reg[8]  ( .CR(1'b1), .D(stage4[8]), .LD(n365), .CP(clock), .Q(
        stage5[8]) );
  FDS2L \stage5_reg[7]  ( .CR(1'b1), .D(stage4[7]), .LD(n365), .CP(clock), .Q(
        stage5[7]) );
  FDS2L \stage5_reg[6]  ( .CR(1'b1), .D(stage4[6]), .LD(n365), .CP(clock), .Q(
        stage5[6]) );
  FDS2L \stage5_reg[5]  ( .CR(1'b1), .D(stage4[5]), .LD(n365), .CP(clock), .Q(
        stage5[5]) );
  FDS2L \stage5_reg[4]  ( .CR(1'b1), .D(stage4[4]), .LD(n365), .CP(clock), .Q(
        stage5[4]) );
  FDS2L \stage5_reg[3]  ( .CR(1'b1), .D(stage4[3]), .LD(n365), .CP(clock), .Q(
        stage5[3]) );
  FDS2L \stage5_reg[2]  ( .CR(1'b1), .D(stage4[2]), .LD(n365), .CP(clock), .Q(
        stage5[2]) );
  FDS2L \stage5_reg[1]  ( .CR(1'b1), .D(stage4[1]), .LD(n365), .CP(clock), .Q(
        stage5[1]) );
  FDS2L \stage5_reg[0]  ( .CR(1'b1), .D(stage4[0]), .LD(n365), .CP(clock), .Q(
        stage5[0]) );
  FDS2L \stage6_reg[16]  ( .CR(1'b1), .D(stage5[16]), .LD(n365), .CP(clock), 
        .Q(stage6[16]) );
  FDS2L \stage6_reg[15]  ( .CR(1'b1), .D(stage5[15]), .LD(n365), .CP(clock), 
        .Q(stage6[15]) );
  FDS2L \stage6_reg[14]  ( .CR(1'b1), .D(stage5[14]), .LD(n365), .CP(clock), 
        .Q(stage6[14]) );
  FDS2L \stage6_reg[13]  ( .CR(1'b1), .D(stage5[13]), .LD(n365), .CP(clock), 
        .Q(stage6[13]) );
  FDS2L \stage6_reg[12]  ( .CR(1'b1), .D(stage5[12]), .LD(n365), .CP(clock), 
        .Q(stage6[12]) );
  FDS2L \stage6_reg[11]  ( .CR(1'b1), .D(stage5[11]), .LD(n365), .CP(clock), 
        .Q(stage6[11]) );
  FDS2L \stage6_reg[10]  ( .CR(1'b1), .D(stage5[10]), .LD(n365), .CP(clock), 
        .Q(stage6[10]) );
  FDS2L \stage6_reg[9]  ( .CR(1'b1), .D(stage5[9]), .LD(n365), .CP(clock), .Q(
        stage6[9]) );
  FDS2L \stage6_reg[8]  ( .CR(1'b1), .D(stage5[8]), .LD(n365), .CP(clock), .Q(
        stage6[8]) );
  FDS2L \stage6_reg[7]  ( .CR(1'b1), .D(stage5[7]), .LD(n365), .CP(clock), .Q(
        stage6[7]) );
  FDS2L \stage6_reg[6]  ( .CR(1'b1), .D(stage5[6]), .LD(n365), .CP(clock), .Q(
        stage6[6]) );
  FDS2L \stage6_reg[5]  ( .CR(1'b1), .D(stage5[5]), .LD(n365), .CP(clock), .Q(
        stage6[5]) );
  FDS2L \stage6_reg[4]  ( .CR(1'b1), .D(stage5[4]), .LD(n365), .CP(clock), .Q(
        stage6[4]) );
  FDS2L \stage6_reg[3]  ( .CR(1'b1), .D(stage5[3]), .LD(n365), .CP(clock), .Q(
        stage6[3]) );
  FDS2L \stage6_reg[2]  ( .CR(1'b1), .D(stage5[2]), .LD(n365), .CP(clock), .Q(
        stage6[2]) );
  FDS2L \stage6_reg[1]  ( .CR(1'b1), .D(stage5[1]), .LD(n365), .CP(clock), .Q(
        stage6[1]) );
  FDS2L \stage6_reg[0]  ( .CR(1'b1), .D(stage5[0]), .LD(n365), .CP(clock), .Q(
        stage6[0]) );
  FD1 \X0_reg[15]  ( .D(N50), .CP(clock), .Q(X0[15]) );
  FD1 \X1_reg[15]  ( .D(N66), .CP(clock), .Q(X1[15]) );
  FDS2L \X0_reg_reg[31]  ( .CR(1'b1), .D(N19), .LD(n365), .CP(clock), .Q(
        X0_reg[31]) );
  FDS2 \X0_reg[14]  ( .CR(X0_reg[31]), .D(n365), .CP(clock), .Q(X0[14]) );
  FDS2L \X0_reg_reg[30]  ( .CR(1'b1), .D(N18), .LD(n365), .CP(clock), .Q(
        X0_reg[30]) );
  FDS2 \X0_reg[13]  ( .CR(X0_reg[30]), .D(n365), .CP(clock), .Q(X0[13]) );
  FDS2L \X0_reg_reg[29]  ( .CR(1'b1), .D(N17), .LD(n365), .CP(clock), .Q(
        X0_reg[29]) );
  FDS2 \X0_reg[12]  ( .CR(X0_reg[29]), .D(n365), .CP(clock), .Q(X0[12]) );
  FDS2L \X0_reg_reg[28]  ( .CR(1'b1), .D(N16), .LD(n365), .CP(clock), .Q(
        X0_reg[28]) );
  FDS2 \X0_reg[11]  ( .CR(X0_reg[28]), .D(n365), .CP(clock), .Q(X0[11]) );
  FDS2L \X0_reg_reg[27]  ( .CR(1'b1), .D(N15), .LD(n365), .CP(clock), .Q(
        X0_reg[27]) );
  FDS2 \X0_reg[10]  ( .CR(X0_reg[27]), .D(n365), .CP(clock), .Q(X0[10]) );
  FDS2L \X0_reg_reg[26]  ( .CR(1'b1), .D(N14), .LD(n365), .CP(clock), .Q(
        X0_reg[26]) );
  FDS2 \X0_reg[9]  ( .CR(X0_reg[26]), .D(n365), .CP(clock), .Q(X0[9]) );
  FDS2L \X0_reg_reg[25]  ( .CR(1'b1), .D(N13), .LD(n365), .CP(clock), .Q(
        X0_reg[25]) );
  FDS2 \X0_reg[8]  ( .CR(X0_reg[25]), .D(n365), .CP(clock), .Q(X0[8]) );
  FDS2L \X0_reg_reg[24]  ( .CR(1'b1), .D(N12), .LD(n365), .CP(clock), .Q(
        X0_reg[24]) );
  FDS2 \X0_reg[7]  ( .CR(X0_reg[24]), .D(n365), .CP(clock), .Q(X0[7]) );
  FDS2L \X0_reg_reg[23]  ( .CR(1'b1), .D(N11), .LD(n365), .CP(clock), .Q(
        X0_reg[23]) );
  FDS2 \X0_reg[6]  ( .CR(X0_reg[23]), .D(n365), .CP(clock), .Q(X0[6]) );
  FDS2L \X0_reg_reg[22]  ( .CR(1'b1), .D(N10), .LD(n365), .CP(clock), .Q(
        X0_reg[22]) );
  FDS2 \X0_reg[5]  ( .CR(X0_reg[22]), .D(n365), .CP(clock), .Q(X0[5]) );
  FDS2L \X0_reg_reg[21]  ( .CR(1'b1), .D(N9), .LD(n365), .CP(clock), .Q(
        X0_reg[21]) );
  FDS2 \X0_reg[4]  ( .CR(X0_reg[21]), .D(n365), .CP(clock), .Q(X0[4]) );
  FDS2L \X0_reg_reg[20]  ( .CR(1'b1), .D(N8), .LD(n365), .CP(clock), .Q(
        X0_reg[20]) );
  FDS2 \X0_reg[3]  ( .CR(X0_reg[20]), .D(n365), .CP(clock), .Q(X0[3]) );
  FDS2L \X0_reg_reg[19]  ( .CR(1'b1), .D(N7), .LD(n365), .CP(clock), .Q(
        X0_reg[19]) );
  FDS2 \X0_reg[2]  ( .CR(X0_reg[19]), .D(n365), .CP(clock), .Q(X0[2]) );
  FDS2L \X0_reg_reg[18]  ( .CR(1'b1), .D(N6), .LD(n365), .CP(clock), .Q(
        X0_reg[18]) );
  FDS2 \X0_reg[1]  ( .CR(X0_reg[18]), .D(n365), .CP(clock), .Q(X0[1]) );
  FDS2L \X0_reg_reg[17]  ( .CR(1'b1), .D(N5), .LD(n365), .CP(clock), .Q(
        X0_reg[17]) );
  FDS2 \X0_reg[0]  ( .CR(X0_reg[17]), .D(n365), .CP(clock), .Q(X0[0]) );
  FDS2L \X1_reg_reg[31]  ( .CR(1'b1), .D(N34), .LD(n365), .CP(clock), .Q(
        X1_reg[31]) );
  FDS2 \X1_reg[14]  ( .CR(X1_reg[31]), .D(n365), .CP(clock), .Q(X1[14]) );
  FDS2L \X1_reg_reg[30]  ( .CR(1'b1), .D(N33), .LD(n365), .CP(clock), .Q(
        X1_reg[30]) );
  FDS2 \X1_reg[13]  ( .CR(X1_reg[30]), .D(n365), .CP(clock), .Q(X1[13]) );
  FDS2L \X1_reg_reg[29]  ( .CR(1'b1), .D(N32), .LD(n365), .CP(clock), .Q(
        X1_reg[29]) );
  FDS2 \X1_reg[12]  ( .CR(X1_reg[29]), .D(n365), .CP(clock), .Q(X1[12]) );
  FDS2L \X1_reg_reg[28]  ( .CR(1'b1), .D(N31), .LD(n365), .CP(clock), .Q(
        X1_reg[28]) );
  FDS2 \X1_reg[11]  ( .CR(X1_reg[28]), .D(n365), .CP(clock), .Q(X1[11]) );
  FDS2L \X1_reg_reg[27]  ( .CR(1'b1), .D(N30), .LD(n365), .CP(clock), .Q(
        X1_reg[27]) );
  FDS2 \X1_reg[10]  ( .CR(X1_reg[27]), .D(n365), .CP(clock), .Q(X1[10]) );
  FDS2L \X1_reg_reg[26]  ( .CR(1'b1), .D(N29), .LD(n365), .CP(clock), .Q(
        X1_reg[26]) );
  FDS2 \X1_reg[9]  ( .CR(X1_reg[26]), .D(n365), .CP(clock), .Q(X1[9]) );
  FDS2L \X1_reg_reg[25]  ( .CR(1'b1), .D(N28), .LD(n365), .CP(clock), .Q(
        X1_reg[25]) );
  FDS2 \X1_reg[8]  ( .CR(X1_reg[25]), .D(n365), .CP(clock), .Q(X1[8]) );
  FDS2L \X1_reg_reg[24]  ( .CR(1'b1), .D(N27), .LD(n365), .CP(clock), .Q(
        X1_reg[24]) );
  FDS2 \X1_reg[7]  ( .CR(X1_reg[24]), .D(n365), .CP(clock), .Q(X1[7]) );
  FDS2L \X1_reg_reg[23]  ( .CR(1'b1), .D(N26), .LD(n365), .CP(clock), .Q(
        X1_reg[23]) );
  FDS2 \X1_reg[6]  ( .CR(X1_reg[23]), .D(n365), .CP(clock), .Q(X1[6]) );
  FDS2L \X1_reg_reg[22]  ( .CR(1'b1), .D(N25), .LD(n365), .CP(clock), .Q(
        X1_reg[22]) );
  FDS2 \X1_reg[5]  ( .CR(X1_reg[22]), .D(n365), .CP(clock), .Q(X1[5]) );
  FDS2L \X1_reg_reg[21]  ( .CR(1'b1), .D(N24), .LD(n365), .CP(clock), .Q(
        X1_reg[21]) );
  FDS2 \X1_reg[4]  ( .CR(X1_reg[21]), .D(n365), .CP(clock), .Q(X1[4]) );
  FDS2L \X1_reg_reg[20]  ( .CR(1'b1), .D(N23), .LD(n365), .CP(clock), .Q(
        X1_reg[20]) );
  FDS2 \X1_reg[3]  ( .CR(X1_reg[20]), .D(n365), .CP(clock), .Q(X1[3]) );
  FDS2L \X1_reg_reg[19]  ( .CR(1'b1), .D(N22), .LD(n365), .CP(clock), .Q(
        X1_reg[19]) );
  FDS2 \X1_reg[2]  ( .CR(X1_reg[19]), .D(n365), .CP(clock), .Q(X1[2]) );
  FDS2L \X1_reg_reg[18]  ( .CR(1'b1), .D(N21), .LD(n365), .CP(clock), .Q(
        X1_reg[18]) );
  FDS2 \X1_reg[1]  ( .CR(X1_reg[18]), .D(n365), .CP(clock), .Q(X1[1]) );
  FDS2L \X1_reg_reg[17]  ( .CR(1'b1), .D(N20), .LD(n365), .CP(clock), .Q(
        X1_reg[17]) );
  FDS2 \X1_reg[0]  ( .CR(X1_reg[17]), .D(n365), .CP(clock), .Q(X1[0]) );
  FDS2L \X01_reg[15]  ( .CR(1'b1), .D(X0[15]), .LD(n365), .CP(clock), .Q(
        X01[15]) );
  FDS2L \X01_reg[14]  ( .CR(1'b1), .D(X0[14]), .LD(n365), .CP(clock), .Q(
        X01[14]) );
  FDS2L \X01_reg[13]  ( .CR(1'b1), .D(X0[13]), .LD(n365), .CP(clock), .Q(
        X01[13]) );
  FDS2L \X01_reg[12]  ( .CR(1'b1), .D(X0[12]), .LD(n365), .CP(clock), .Q(
        X01[12]) );
  FDS2L \X01_reg[11]  ( .CR(1'b1), .D(X0[11]), .LD(n365), .CP(clock), .Q(
        X01[11]) );
  FDS2L \X01_reg[10]  ( .CR(1'b1), .D(X0[10]), .LD(n365), .CP(clock), .Q(
        X01[10]) );
  FDS2L \X01_reg[9]  ( .CR(1'b1), .D(X0[9]), .LD(n365), .CP(clock), .Q(X01[9])
         );
  FDS2L \X01_reg[8]  ( .CR(1'b1), .D(X0[8]), .LD(n365), .CP(clock), .Q(X01[8])
         );
  FDS2L \X01_reg[7]  ( .CR(1'b1), .D(X0[7]), .LD(n365), .CP(clock), .Q(X01[7])
         );
  FDS2L \X01_reg[6]  ( .CR(1'b1), .D(X0[6]), .LD(n365), .CP(clock), .Q(X01[6])
         );
  FDS2L \X01_reg[5]  ( .CR(1'b1), .D(X0[5]), .LD(n365), .CP(clock), .Q(X01[5])
         );
  FDS2L \X01_reg[4]  ( .CR(1'b1), .D(X0[4]), .LD(n365), .CP(clock), .Q(X01[4])
         );
  FDS2L \X01_reg[3]  ( .CR(1'b1), .D(X0[3]), .LD(n365), .CP(clock), .Q(X01[3])
         );
  FDS2L \X01_reg[2]  ( .CR(1'b1), .D(X0[2]), .LD(n365), .CP(clock), .Q(X01[2])
         );
  FDS2L \X01_reg[1]  ( .CR(1'b1), .D(X0[1]), .LD(n365), .CP(clock), .Q(X01[1])
         );
  FDS2L \X01_reg[0]  ( .CR(1'b1), .D(X0[0]), .LD(n365), .CP(clock), .Q(X01[0])
         );
  FDS2L \X11_reg[15]  ( .CR(1'b1), .D(X1[15]), .LD(n365), .CP(clock), .Q(
        X11[15]) );
  FDS2L \X11_reg[14]  ( .CR(1'b1), .D(X1[14]), .LD(n365), .CP(clock), .Q(
        X11[14]) );
  FDS2L \X11_reg[13]  ( .CR(1'b1), .D(X1[13]), .LD(n365), .CP(clock), .Q(
        X11[13]) );
  FDS2L \X11_reg[12]  ( .CR(1'b1), .D(X1[12]), .LD(n365), .CP(clock), .Q(
        X11[12]) );
  FDS2L \X11_reg[11]  ( .CR(1'b1), .D(X1[11]), .LD(n365), .CP(clock), .Q(
        X11[11]) );
  FDS2L \X11_reg[10]  ( .CR(1'b1), .D(X1[10]), .LD(n365), .CP(clock), .Q(
        X11[10]) );
  FDS2L \X11_reg[9]  ( .CR(1'b1), .D(X1[9]), .LD(n365), .CP(clock), .Q(X11[9])
         );
  FDS2L \X11_reg[8]  ( .CR(1'b1), .D(X1[8]), .LD(n365), .CP(clock), .Q(X11[8])
         );
  FDS2L \X11_reg[7]  ( .CR(1'b1), .D(X1[7]), .LD(n365), .CP(clock), .Q(X11[7])
         );
  FDS2L \X11_reg[6]  ( .CR(1'b1), .D(X1[6]), .LD(n365), .CP(clock), .Q(X11[6])
         );
  FDS2L \X11_reg[5]  ( .CR(1'b1), .D(X1[5]), .LD(n365), .CP(clock), .Q(X11[5])
         );
  FDS2L \X11_reg[4]  ( .CR(1'b1), .D(X1[4]), .LD(n365), .CP(clock), .Q(X11[4])
         );
  FDS2L \X11_reg[3]  ( .CR(1'b1), .D(X1[3]), .LD(n365), .CP(clock), .Q(X11[3])
         );
  FDS2L \X11_reg[2]  ( .CR(1'b1), .D(X1[2]), .LD(n365), .CP(clock), .Q(X11[2])
         );
  FDS2L \X11_reg[1]  ( .CR(1'b1), .D(X1[1]), .LD(n365), .CP(clock), .Q(X11[1])
         );
  FDS2L \X11_reg[0]  ( .CR(1'b1), .D(X1[0]), .LD(n365), .CP(clock), .Q(X11[0])
         );
  MUX21H U317 ( .A(Angle[3]), .B(taus_out_0[3]), .S(n365), .Z(n350) );
  MUX21H U318 ( .A(Angle[7]), .B(taus_out_0[7]), .S(n365), .Z(n351) );
  MUX21H U319 ( .A(Angle[11]), .B(taus_out_0[11]), .S(n365), .Z(n352) );
  MUX21H U320 ( .A(Angle[15]), .B(taus_out_0[15]), .S(n365), .Z(n353) );
  MUX21H U321 ( .A(Angle[4]), .B(taus_out_0[4]), .S(n365), .Z(n354) );
  MUX21H U322 ( .A(Angle[8]), .B(taus_out_0[8]), .S(n365), .Z(n355) );
  MUX21H U323 ( .A(Angle[12]), .B(taus_out_0[12]), .S(n365), .Z(n356) );
  MUX21H U324 ( .A(Angle[5]), .B(taus_out_0[5]), .S(n365), .Z(n357) );
  MUX21H U325 ( .A(Angle[9]), .B(taus_out_0[9]), .S(n365), .Z(n358) );
  MUX21H U326 ( .A(Angle[13]), .B(taus_out_0[13]), .S(n365), .Z(n359) );
  MUX21H U327 ( .A(Angle[6]), .B(taus_out_0[6]), .S(n365), .Z(n360) );
  MUX21H U328 ( .A(Angle[10]), .B(taus_out_0[10]), .S(n365), .Z(n361) );
  MUX21H U329 ( .A(Angle[14]), .B(taus_out_0[14]), .S(n365), .Z(n362) );
  MUX21H U330 ( .A(Angle[2]), .B(taus_out_0[2]), .S(n365), .Z(n363) );
  MUX21H U331 ( .A(Angle[1]), .B(taus_out_0[1]), .S(n365), .Z(n364) );
  AN2 U332 ( .A(cos_out[15]), .B(n365), .Z(N66) );
  AN2 U333 ( .A(sin_out[15]), .B(n365), .Z(N50) );
  IV U334 ( .A(reset), .Z(n365) );
endmodule

