 //Awgn using box_muller_method
//Rahul Umrania
//W1114663

//Top Module//

module top_module(clock, reset, X0_output, X1_output, valid);
input clock;
input reset;

output reg [15:0] X0_output;
output reg[15:0] X1_output;
output reg valid;
wire  [15:0] cos_out;
wire  [15:0] sin_out;

localparam VALUE = 32000/1.647; //Xin for Cordic
// tausworthe generator 
wire [31:0] taus_out_0;
wire [31:0] taus_out_1;
reg [15:0] Angle, X01, X11,X0, X1;

//logarithm out block
reg [30:0] LogOut2;
wire [30:0] logarith_out;
reg [47:0] LogIn;
// square out 
wire [16:0] sqrt_out;
reg [16:0] stage0, stage1, stage2, stage3, stage4, stage5, stage6, sqrtOut;
reg valid0, valid1, valid2, valid3, valid4, valid5, valid6, valid7, valid8, valid9, valid10, valid11, valid12, valid13, valid14, valid15;

// sin/cos
wire [15:0] x_out;
wire [15:0] y_out;

reg [31:0] X0_reg, X1_reg;

	always @(posedge clock) begin
		
		valid0 <= !reset;
		valid1 <= valid0;
		valid2 <= valid1;
		valid3 <= valid2;
		valid4 <= valid3;
		valid5 <= valid4;
		valid6 <= valid5;
		valid7 <= valid6;
		valid8 <= valid7;
		valid9 <= valid8;
		valid10 <= valid9;
		valid11 <= valid10;
		valid12 <= valid11;
		valid13 <= valid12;
		valid14 <= valid13;
		valid15 <= valid14;
		valid <= valid15;
			
	
		if(!reset) begin

			LogIn <= {taus_out_1[31:0], taus_out_0[31:16]};
			Angle <= taus_out_0[15:0];

			stage0 <= sqrt_out;
			stage1 <= stage0;
			stage2 <= stage1;
			stage3 <= stage2;
			stage4 <= stage3;
			stage5 <= stage4;
			stage6 <= stage5;
			sqrtOut <= stage6;

			LogOut2 <= logarith_out;
		
			X0[15] <= sin_out[15];
			X1[15] <= cos_out[15];
			
			X0_reg <= sin_out[14:0] * sqrtOut[16:0];
			X1_reg <= cos_out[14:0] * sqrtOut[16:0];
			
			X0[14:11] <= X0_reg[31:28];
			X0[10:0] <= X0_reg[27:17];

			X1[14:11] <= X1_reg[31:28];
			X1[10:0] <= X1_reg[27:17];
			
		X01 <= X0;
		X11 <= X1;

		X0_output <= X01;
		X1_output <= X11;

		end
			
		else begin
			valid <= 1'b0;
			valid0 <= 1'b0;
			valid1 <= 1'b0;
			valid2 <= 1'b0;
			valid3 <= 1'b0;
			valid4 <= 1'b0;
			valid5 <= 1'b0;
			valid6 <= 1'b0;
			valid7 <= 1'b0;
			valid8 <= 1'b0;
			valid9 <= 1'b0;
			valid10 <= 1'b0;
			valid11 <= 1'b0;
			valid12 <= 1'b0;
			valid13 <= 1'b0;
			valid14 <= 1'b0;
			valid15 <= 1'b0;

			X0 <= 15'b0;
			X1 <= 15'b0;
		end

	
	end
	

tausworthe taus_gen (clock, reset, taus_out_0);
tausworthe taus_gen1(clock, reset, taus_out_1);
CORDIC codic_sin_cos (clock, Angle, VALUE, 16'b0, cos_out, sin_out);
Poly_Logarithm login(clock, reset, LogIn , logarith_out);
Poly_sqrt sqrt1 (clock, reset, logarith_out, sqrt_out);

endmodule





module tausworthe (clock, re_set, tausout);

//***Define the Parameter_width*****//
	parameter width = 32;
	
//***Define the inputs*********//
	input clock;
	input re_set;
	
//***Define the outputs********//
	output [width-1:0] tausout ;
	
	reg [width-1:0] Seed_0;
	reg [width-1:0] Seed_1;
	reg [width-1:0] Seed_2;
	reg [width-1:0] b;
//***Assigning tausout********//
	assign tausout = Seed_0 ^ Seed_1 ^ Seed_2;
	always @ (posedge clock ) begin
		if(!re_set) begin
	
			b = ((( Seed_0 << 13) ^ Seed_0) >> 19);

			Seed_0 = ((( Seed_0 & 32'hFFFFFFFE) << 12 ) ^ b);

			b = ((( Seed_1 << 2) ^ Seed_1) >> 25);

			Seed_1 = ((( Seed_1 & 32'hFFFF_FFF8) << 4 ) ^ b);

			b = ((( Seed_2 << 3) ^ Seed_2) >> 11);
	
			Seed_2 = ((( Seed_2 & 32'hFFFF_FFF0) << 17 ) ^ b);
		end
		else begin
			Seed_0 = 4;
			Seed_1 = 5;
			Seed_2 = 7;
		end
	end
endmodule

// module Cordic 
// NOTE: 1. Input angle is a modulo of 2*PI scaled to fit in a 32bit register. The user must translate
//          this angle to a value from 0 - (2^32-1).  0 deg = 32'h0, 359.9999... = 32'hFF_FF_FF_FF
//          To translate from degrees to a 32 bit value, multiply 2^32 by the angle (in degrees),
//          then divide by 360
//       2. Size of cos_out, sin_out is 1 bit larger due to a system gain of 1.647 (which is < 2)
module CORDIC (clock, angle, Xin, Yin, cos_out, sin_out);
   
   parameter XY_SZ = 16;   // width of input and output data
   
   localparam STG = XY_SZ; // same as bit width of X and Y
   
   input                      clock;
   // angle is a signed value in the range of -PI to +PI that must be represented as a 32 bit signed number
   input         [15:0] angle;
   input      [XY_SZ-1:0] Xin;
   input      [XY_SZ-1:0] Yin;
   output      [XY_SZ-1:0] cos_out;
   output      [XY_SZ-1:0] sin_out;
   
   //------------------------------------------------------------------------------
   //                             arctan table
   //------------------------------------------------------------------------------
   
   // Note: The atan_table was chosen to be 31 bits wide giving resolution up to atan(2^-30)
   wire  [31:0] atan_table [0:30];
   
   // upper 2 bits = 2'b00 which represents 0 - PI/2 range
   // upper 2 bits = 2'b01 which represents PI/2 to PI range
   // upper 2 bits = 2'b10 which represents PI to 3*PI/2 range (i.e. -PI/2 to -PI)
   // upper 2 bits = 2'b11 which represents 3*PI/2 to 2*PI range (i.e. 0 to -PI/2)
   // The upper 2 bits therefore tell us which quadrant we are in.
   assign atan_table[00] = 32'b00100000000000000000000000000000; // 45.000 degrees -> atan(2^0)
   assign atan_table[01] = 32'b00010010111001000000010100011101; // 26.565 degrees -> atan(2^-1)
   assign atan_table[02] = 32'b00001001111110110011100001011011; // 14.036 degrees -> atan(2^-2)
   assign atan_table[03] = 32'b00000101000100010001000111010100; // atan(2^-3)
   assign atan_table[04] = 32'b00000010100010110000110101000011;
   assign atan_table[05] = 32'b00000001010001011101011111100001;
   assign atan_table[06] = 32'b00000000101000101111011000011110;
   assign atan_table[07] = 32'b00000000010100010111110001010101;
   assign atan_table[08] = 32'b00000000001010001011111001010011;
   assign atan_table[09] = 32'b00000000000101000101111100101110;
   assign atan_table[10] = 32'b00000000000010100010111110011000;
   assign atan_table[11] = 32'b00000000000001010001011111001100;
   assign atan_table[12] = 32'b00000000000000101000101111100110;
   assign atan_table[13] = 32'b00000000000000010100010111110011;
   assign atan_table[14] = 32'b00000000000000001010001011111001;
   assign atan_table[15] = 32'b00000000000000000101000101111101;
   assign atan_table[16] = 32'b00000000000000000010100010111110;
   assign atan_table[17] = 32'b00000000000000000001010001011111;
   assign atan_table[18] = 32'b00000000000000000000101000101111;
   assign atan_table[19] = 32'b00000000000000000000010100011000;
   assign atan_table[20] = 32'b00000000000000000000001010001100;
   assign atan_table[21] = 32'b00000000000000000000000101000110;
   assign atan_table[22] = 32'b00000000000000000000000010100011;
   assign atan_table[23] = 32'b00000000000000000000000001010001;
   assign atan_table[24] = 32'b00000000000000000000000000101000;
   assign atan_table[25] = 32'b00000000000000000000000000010100;
   assign atan_table[26] = 32'b00000000000000000000000000001010;
   assign atan_table[27] = 32'b00000000000000000000000000000101;
   assign atan_table[28] = 32'b00000000000000000000000000000010;
   assign atan_table[29] = 32'b00000000000000000000000000000001; // atan(2^-29)
   assign atan_table[30] = 32'b00000000000000000000000000000000;
   
   //------------------------------------------------------------------------------
   //                              registers
   //------------------------------------------------------------------------------
   
   //stage outputs
   reg  [XY_SZ:0] X [0:STG-1];
   reg  [XY_SZ:0] Y [0:STG-1];
   reg     [31:0] Z [0:STG-1]; // 32bit
   
   //------------------------------------------------------------------------------
   //                               stage 0
   //------------------------------------------------------------------------------
   wire                 [1:0] quadrant;
   assign   quadrant = angle[15:14];
   
   always @(posedge clock)
   begin // make sure the rotation angle is in the -pi/2 to pi/2 range.  If not then pre-rotate
      case (quadrant)
         2'b00,
         2'b11:   // no pre-rotation needed for these quadrants
         begin    // X[n], Y[n] is 1 bit larger than Xin, Yin, but Verilog handles the assignments properly
            X[0] <= Xin;
            Y[0] <= Yin;
            Z[0] <= angle;
         end
         
         2'b01:
         begin
            X[0] <= -Yin;
            Y[0] <= Xin;
            Z[0] <= {2'b00,angle[13:0]}; // subtract pi/2 from angle for this quadrant
         end
         
         2'b10:
         begin
            X[0] <= Yin;
            Y[0] <= -Xin;
            Z[0] <= {2'b11,angle[13:0]}; // add pi/2 to angle for this quadrant
         end
         
      endcase
   end
   
   //------------------------------------------------------------------------------
   //                           generate stages 1 to STG-1
   //------------------------------------------------------------------------------
   genvar i;

   generate
   for (i=0; i < (STG-1); i=i+1)
   begin: XYZ
      wire                   Z_sign;
      wire  [XY_SZ:0] X_shr, Y_shr; 
   
      assign X_shr = X[i] >>> i; // signed shift right
      assign Y_shr = Y[i] >>> i;
   
      //the sign of the current rotation angle
      assign Z_sign = Z[i][15]; // Z_sign = 1 if Z[i] < 0
   
      always @(posedge clock)
      begin
         // add/subtract shifted data
         X[i+1] <= Z_sign ? X[i] + Y_shr         : X[i] - Y_shr;
         Y[i+1] <= Z_sign ? Y[i] - X_shr         : Y[i] + X_shr;
         Z[i+1] <= Z_sign ? Z[i] + atan_table[i] : Z[i] - atan_table[i];
      end
   end
   endgenerate
   
   
   //------------------------------------------------------------------------------
   //                                 output
   //------------------------------------------------------------------------------
   assign cos_out = X[STG-1];
   assign sin_out = Y[STG-1];

endmodule



/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module Poly_Logarithm(clock, reset, input_log, output_log);
input clock; 
input reset; 
input [47:0] input_log;
output reg [30:0] output_log;


reg [21:0] coeff_log1[256];
reg [12:0] coeff_log0[256];
reg [29:0] coeff_log2[256];
reg [95:0] input_logsquare;
reg [125:0] num1;
reg [69:0] num2;
reg [26:0] num3;

reg [23:0] Fraction_bit;
reg [6:0] Integer_bit;
reg [29:0] Log;

reg [47:0] input_log2;
reg [125:0] num1_1;
reg [69:0] num2_1;
reg [26:0] num3_1;
reg [22:0] Log_P;

always @(posedge clock)
begin
	if(!reset)
	begin

	
		input_logsquare <= input_log * input_log; //square the input
		input_log2 <= input_log;	 
		
		num1 <= input_log * coeff_log2[input_log2[47:40]];
		num2 <= input_log2 * coeff_log1[input_log2[47:40]];
		num3 <= { coeff_log0[input_log2[47:40]], 14'b00000000_000000 };
		
		num1_1 <= num1; // store num1 
		num2_1 <= num2; // store num2 
		num3_1 <= num3; // store num3 

		Fraction_bit <= num1[111:89] - num2[60:38] + num3 [23:1];

	
		Integer_bit <=  num1_1[118:112] - num2_1[67:61] + num3_1 [26:24] + Fraction_bit[23];
		Log_P[22:0] <= Fraction_bit[22:0];

	
		Log[22:0] <= Log_P[22:0];
		Log[29:23] <= Integer_bit[6:0];

		output_log <= Log * 2;

	end

	else begin

		//output_log <= 31'b0;

		//coeff_log2 Coefficient Table

		coeff_log2[0] <= 30'b111111111111111111111111111111;
		coeff_log2[1] <= 30'b111011110010100011100010001111;
		coeff_log2[2] <= 30'b010100110101110010110001110101;
		coeff_log2[3] <= 30'b001010100010101011001001011011;
		coeff_log2[4] <= 30'b000110010110101101001111011101;
		coeff_log2[5] <= 30'b000100001111110001101111110100;
		coeff_log2[6] <= 30'b000011000010011000111000010010;
		coeff_log2[7] <= 30'b000010010001111010100010101111;
		coeff_log2[8] <= 30'b000001110001100011011001111100;
		coeff_log2[9] <= 30'b000001011010111000001110000011;
		coeff_log2[10] <= 30'b000001001010011000000101111001;
		coeff_log2[11] <= 30'b000000111101111111100110010010;
		coeff_log2[12] <= 30'b000000110100011101110000010101;
		coeff_log2[13] <= 30'b000000101100111110011100110111;
		coeff_log2[14] <= 30'b000000100110111110111010101110;
		coeff_log2[15] <= 30'b000000100010000111001111001110;
		coeff_log2[16] <= 30'b000000011110000110100001010100;
		coeff_log2[17] <= 30'b000000011010110000100011111111;
		coeff_log2[18] <= 30'b000000010111111100010111100010;
		coeff_log2[19] <= 30'b000000010101100011001100000011;
		coeff_log2[20] <= 30'b000000010011011111111000011011;
		coeff_log2[21] <= 30'b000000010001101110011110010000;
		coeff_log2[22] <= 30'b000000010000001011110110011101;
		coeff_log2[23] <= 30'b000000001110110101100011010101;
		coeff_log2[24] <= 30'b000000001101101001100110110010;
		coeff_log2[25] <= 30'b000000001100100110011010111001;
		coeff_log2[26] <= 30'b000000001011101010101100101001;
		coeff_log2[27] <= 30'b000000001010110101010111110100;
		coeff_log2[28] <= 30'b000000001010000101100011111100;
		coeff_log2[29] <= 30'b000000001001011010100010000000;
		coeff_log2[30] <= 30'b000000001000110011101010100001;
		coeff_log2[31] <= 30'b000000001000010000011100001011;
		coeff_log2[32] <= 30'b000000000111110000011010110000;
		coeff_log2[33] <= 30'b000000000111010011001110000111;
		coeff_log2[34] <= 30'b000000000110111000100001101000;
		coeff_log2[35] <= 30'b000000000110100000000011011111;
		coeff_log2[36] <= 30'b000000000110001001100100010101;
		coeff_log2[37] <= 30'b000000000101110100110110110000;
		coeff_log2[38] <= 30'b000000000101100001101111001001;
		coeff_log2[39] <= 30'b000000000101010000000011010010;
		coeff_log2[40] <= 30'b000000000100111111101010010000;
		coeff_log2[41] <= 30'b000000000100110000011100001000;
		coeff_log2[42] <= 30'b000000000100100010010001111101;
		coeff_log2[43] <= 30'b000000000100010101000101100100;
		coeff_log2[44] <= 30'b000000000100001000110001011110;
		coeff_log2[45] <= 30'b000000000011111101010000110000;
		coeff_log2[46] <= 30'b000000000011110010011111000100;
		coeff_log2[47] <= 30'b000000000011101000011000011111;
		coeff_log2[48] <= 30'b000000000011011110111001011110;
		coeff_log2[49] <= 30'b000000000011010101111110111001;
		coeff_log2[50] <= 30'b000000000011001101100101110111;
		coeff_log2[51] <= 30'b000000000011000101101011110101;
		coeff_log2[52] <= 30'b000000000010111110001110011011;
		coeff_log2[53] <= 30'b000000000010110111001011100010;
		coeff_log2[54] <= 30'b000000000010110000100001010000;
		coeff_log2[55] <= 30'b000000000010101010001101110011;
		coeff_log2[56] <= 30'b000000000010100100001111100101;
		coeff_log2[57] <= 30'b000000000010011110100101001000;
		coeff_log2[58] <= 30'b000000000010011001001101000110;
		coeff_log2[59] <= 30'b000000000010010100000110010001;
		coeff_log2[60] <= 30'b000000000010001111001111100001;
		coeff_log2[61] <= 30'b000000000010001010100111110100;
		coeff_log2[62] <= 30'b000000000010000110001110001011;
		coeff_log2[63] <= 30'b000000000010000010000001101111;
		coeff_log2[64] <= 30'b000000000001111110000001101100;
		coeff_log2[65] <= 30'b000000000001111010001101010010;
		coeff_log2[66] <= 30'b000000000001110110100011110101;
		coeff_log2[67] <= 30'b000000000001110011000100101010;
		coeff_log2[68] <= 30'b000000000001101111101111001101;
		coeff_log2[69] <= 30'b000000000001101100100010111000;
		coeff_log2[70] <= 30'b000000000001101001011111001101;
		coeff_log2[71] <= 30'b000000000001100110100011101011;
		coeff_log2[72] <= 30'b000000000001100011101111110110;
		coeff_log2[73] <= 30'b000000000001100001000011010100;
		coeff_log2[74] <= 30'b000000000001011110011101101100;
		coeff_log2[75] <= 30'b000000000001011011111110100110;
		coeff_log2[76] <= 30'b000000000001011001100101101101;
		coeff_log2[77] <= 30'b000000000001010111010010101100;
		coeff_log2[78] <= 30'b000000000001010101000101010000;
		coeff_log2[79] <= 30'b000000000001010010111101001000;
		coeff_log2[80] <= 30'b000000000001010000111010000011;
		coeff_log2[81] <= 30'b000000000001001110111011110000;
		coeff_log2[82] <= 30'b000000000001001101000010000001;
		coeff_log2[83] <= 30'b000000000001001011001100101001;
		coeff_log2[84] <= 30'b000000000001001001011011011010;
		coeff_log2[85] <= 30'b000000000001000111101110001000;
		coeff_log2[86] <= 30'b000000000001000110000100100111;
		coeff_log2[87] <= 30'b000000000001000100011110101100;
		coeff_log2[88] <= 30'b000000000001000010111100001101;
		coeff_log2[89] <= 30'b000000000001000001011101000000;
		coeff_log2[90] <= 30'b000000000001000000000000111011;
		coeff_log2[91] <= 30'b000000000000111110100111110111;
		coeff_log2[92] <= 30'b000000000000111101010001101011;
		coeff_log2[93] <= 30'b000000000000111011111110001111;
		coeff_log2[94] <= 30'b000000000000111010101101011100;
		coeff_log2[95] <= 30'b000000000000111001011111001010;
		coeff_log2[96] <= 30'b000000000000111000010011010011;
		coeff_log2[97] <= 30'b000000000000110111001001110001;
		coeff_log2[98] <= 30'b000000000000110110000010011101;
		coeff_log2[99] <= 30'b000000000000110100111101010010;
		coeff_log2[100] <= 30'b000000000000110011111010001011;
		coeff_log2[101] <= 30'b000000000000110010111001000010;
		coeff_log2[102] <= 30'b000000000000110001111001110011;
		coeff_log2[103] <= 30'b000000000000110000111100011000;
		coeff_log2[104] <= 30'b000000000000110000000000101101;
		coeff_log2[105] <= 30'b000000000000101111000110101111;
		coeff_log2[106] <= 30'b000000000000101110001110011001;
		coeff_log2[107] <= 30'b000000000000101101010111100110;
		coeff_log2[108] <= 30'b000000000000101100100010010101;
		coeff_log2[109] <= 30'b000000000000101011101110100000;
		coeff_log2[110] <= 30'b000000000000101010111100000101;
		coeff_log2[111] <= 30'b000000000000101010001011000000;
		coeff_log2[112] <= 30'b000000000000101001011011001111;
		coeff_log2[113] <= 30'b000000000000101000101100101110;
		coeff_log2[114] <= 30'b000000000000100111111111011011;
		coeff_log2[115] <= 30'b000000000000100111010011010011;
		coeff_log2[116] <= 30'b000000000000100110101000010011;
		coeff_log2[117] <= 30'b000000000000100101111110011010;
		coeff_log2[118] <= 30'b000000000000100101010101100011;
		coeff_log2[119] <= 30'b000000000000100100101101101111;
		coeff_log2[120] <= 30'b000000000000100100000110111001;
		coeff_log2[121] <= 30'b000000000000100011100001000000;
		coeff_log2[122] <= 30'b000000000000100010111100000011;
		coeff_log2[123] <= 30'b000000000000100010010111111111;
		coeff_log2[124] <= 30'b000000000000100001110100110010;
		coeff_log2[125] <= 30'b000000000000100001010010011011;
		coeff_log2[126] <= 30'b000000000000100000110000111000;
		coeff_log2[127] <= 30'b000000000000100000010000000111;
		coeff_log2[128] <= 30'b000000000000011111110000000111;
		coeff_log2[129] <= 30'b000000000000011111010000110110;
		coeff_log2[130] <= 30'b000000000000011110110010010011;
		coeff_log2[131] <= 30'b000000000000011110010100011100;
		coeff_log2[132] <= 30'b000000000000011101110111010001;
		coeff_log2[133] <= 30'b000000000000011101011010101111;
		coeff_log2[134] <= 30'b000000000000011100111110110110;
		coeff_log2[135] <= 30'b000000000000011100100011100100;
		coeff_log2[136] <= 30'b000000000000011100001000111001;
		coeff_log2[137] <= 30'b000000000000011011101110110011;
		coeff_log2[138] <= 30'b000000000000011011010101010000;
		coeff_log2[139] <= 30'b000000000000011010111100010001;
		coeff_log2[140] <= 30'b000000000000011010100011110100;
		coeff_log2[141] <= 30'b000000000000011010001011110111;
		coeff_log2[142] <= 30'b000000000000011001110100011011;
		coeff_log2[143] <= 30'b000000000000011001011101011111;
		coeff_log2[144] <= 30'b000000000000011001000111000000;
		coeff_log2[145] <= 30'b000000000000011000110000111111;
		coeff_log2[146] <= 30'b000000000000011000011011011011;
		coeff_log2[147] <= 30'b000000000000011000000110010011;
		coeff_log2[148] <= 30'b000000000000010111110001100110;
		coeff_log2[149] <= 30'b000000000000010111011101010100;
		coeff_log2[150] <= 30'b000000000000010111001001011011;
		coeff_log2[151] <= 30'b000000000000010110110101111100;
		coeff_log2[152] <= 30'b000000000000010110100010110100;
		coeff_log2[153] <= 30'b000000000000010110010000000101;
		coeff_log2[154] <= 30'b000000000000010101111101101101;
		coeff_log2[155] <= 30'b000000000000010101101011101100;
		coeff_log2[156] <= 30'b000000000000010101011010000001;
		coeff_log2[157] <= 30'b000000000000010101001000101011;
		coeff_log2[158] <= 30'b000000000000010100110111101010;
		coeff_log2[159] <= 30'b000000000000010100100110111101;
		coeff_log2[160] <= 30'b000000000000010100010110100101;
		coeff_log2[161] <= 30'b000000000000010100000110011111;
		coeff_log2[162] <= 30'b000000000000010011110110101101;
		coeff_log2[163] <= 30'b000000000000010011100111001101;
		coeff_log2[164] <= 30'b000000000000010011011000000000;
		coeff_log2[165] <= 30'b000000000000010011001001000100;
		coeff_log2[166] <= 30'b000000000000010010111010011001;
		coeff_log2[167] <= 30'b000000000000010010101011111110;
		coeff_log2[168] <= 30'b000000000000010010011101110101;
		coeff_log2[169] <= 30'b000000000000010010001111111011;
		coeff_log2[170] <= 30'b000000000000010010000010010000;
		coeff_log2[171] <= 30'b000000000000010001110100110110;
		coeff_log2[172] <= 30'b000000000000010001100111101001;
		coeff_log2[173] <= 30'b000000000000010001011010101100;
		coeff_log2[174] <= 30'b000000000000010001001101111101;
		coeff_log2[175] <= 30'b000000000000010001000001011011;
		coeff_log2[176] <= 30'b000000000000010000110101000111;
		coeff_log2[177] <= 30'b000000000000010000101001000001;
		coeff_log2[178] <= 30'b000000000000010000011101000111;
		coeff_log2[179] <= 30'b000000000000010000010001011010;
		coeff_log2[180] <= 30'b000000000000010000000101111010;
		coeff_log2[181] <= 30'b000000000000001111111010100110;
		coeff_log2[182] <= 30'b000000000000001111101111011101;
		coeff_log2[183] <= 30'b000000000000001111100100100000;
		coeff_log2[184] <= 30'b000000000000001111011001101111;
		coeff_log2[185] <= 30'b000000000000001111001111001000;
		coeff_log2[186] <= 30'b000000000000001111000100101101;
		coeff_log2[187] <= 30'b000000000000001110111010011100;
		coeff_log2[188] <= 30'b000000000000001110110000010110;
		coeff_log2[189] <= 30'b000000000000001110100110011010;
		coeff_log2[190] <= 30'b000000000000001110011100100111;
		coeff_log2[191] <= 30'b000000000000001110010010111111;
		coeff_log2[192] <= 30'b000000000000001110001001100000;
		coeff_log2[193] <= 30'b000000000000001110000000001011;
		coeff_log2[194] <= 30'b000000000000001101110110111110;
		coeff_log2[195] <= 30'b000000000000001101101101111011;
		coeff_log2[196] <= 30'b000000000000001101100101000001;
		coeff_log2[197] <= 30'b000000000000001101011100001111;
		coeff_log2[198] <= 30'b000000000000001101010011100110;
		coeff_log2[199] <= 30'b000000000000001101001011000101;
		coeff_log2[200] <= 30'b000000000000001101000010101100;
		coeff_log2[201] <= 30'b000000000000001100111010011011;
		coeff_log2[202] <= 30'b000000000000001100110010010010;
		coeff_log2[203] <= 30'b000000000000001100101010010000;
		coeff_log2[204] <= 30'b000000000000001100100010010110;
		coeff_log2[205] <= 30'b000000000000001100011010100100;
		coeff_log2[206] <= 30'b000000000000001100010010111001;
		coeff_log2[207] <= 30'b000000000000001100001011010100;
		coeff_log2[208] <= 30'b000000000000001100000011110111;
		coeff_log2[209] <= 30'b000000000000001011111100100001;
		coeff_log2[210] <= 30'b000000000000001011110101010001;
		coeff_log2[211] <= 30'b000000000000001011101110001000;
		coeff_log2[212] <= 30'b000000000000001011100111000101;
		coeff_log2[213] <= 30'b000000000000001011100000001000;
		coeff_log2[214] <= 30'b000000000000001011011001010010;
		coeff_log2[215] <= 30'b000000000000001011010010100010;
		coeff_log2[216] <= 30'b000000000000001011001011111000;
		coeff_log2[217] <= 30'b000000000000001011000101010011;
		coeff_log2[218] <= 30'b000000000000001010111110110101;
		coeff_log2[219] <= 30'b000000000000001010111000011100;
		coeff_log2[220] <= 30'b000000000000001010110010001001;
		coeff_log2[221] <= 30'b000000000000001010101011111011;
		coeff_log2[222] <= 30'b000000000000001010100101110010;
		coeff_log2[223] <= 30'b000000000000001010011111101111;
		coeff_log2[224] <= 30'b000000000000001010011001110001;
		coeff_log2[225] <= 30'b000000000000001010010011111000;
		coeff_log2[226] <= 30'b000000000000001010001110000100;
		coeff_log2[227] <= 30'b000000000000001010001000010100;
		coeff_log2[228] <= 30'b000000000000001010000010101010;
		coeff_log2[229] <= 30'b000000000000001001111101000100;
		coeff_log2[230] <= 30'b000000000000001001110111100011;
		coeff_log2[231] <= 30'b000000000000001001110010000111;
		coeff_log2[232] <= 30'b000000000000001001101100101111;
		coeff_log2[233] <= 30'b000000000000001001100111011011;
		coeff_log2[234] <= 30'b000000000000001001100010001100;
		coeff_log2[235] <= 30'b000000000000001001011101000001;
		coeff_log2[236] <= 30'b000000000000001001010111111010;
		coeff_log2[237] <= 30'b000000000000001001010010111000;
		coeff_log2[238] <= 30'b000000000000001001001101111001;
		coeff_log2[239] <= 30'b000000000000001001001000111111;
		coeff_log2[240] <= 30'b000000000000001001000100001000;
		coeff_log2[241] <= 30'b000000000000001000111111010101;
		coeff_log2[242] <= 30'b000000000000001000111010100110;
		coeff_log2[243] <= 30'b000000000000001000110101111011;
		coeff_log2[244] <= 30'b000000000000001000110001010011;
		coeff_log2[245] <= 30'b000000000000001000101100101111;
		coeff_log2[246] <= 30'b000000000000001000101000001110;
		coeff_log2[247] <= 30'b000000000000001000100011110001;
		coeff_log2[248] <= 30'b000000000000001000011111011000;
		coeff_log2[249] <= 30'b000000000000001000011011000010;
		coeff_log2[250] <= 30'b000000000000001000010110101111;
		coeff_log2[251] <= 30'b000000000000001000010010011111;
		coeff_log2[252] <= 30'b000000000000001000001110010011;
		coeff_log2[253] <= 30'b000000000000001000001010001010;
		coeff_log2[254] <= 30'b000000000000001000000110000011;
		coeff_log2[255] <= 30'b000000000000001000000010000000;


		// Coeff_log1 Table

		coeff_log1[0] <= 22'b1111111111111111111111;
		coeff_log1[1] <= 22'b1011000100000100110111;
		coeff_log1[2] <= 22'b0110011110111000010000;
		coeff_log1[3] <= 22'b0100100110011110011011;
		coeff_log1[4] <= 22'b0011100100011100101001;
		coeff_log1[5] <= 22'b0010111010101010110110;
		coeff_log1[6] <= 22'b0010011101110101010110;
		coeff_log1[7] <= 22'b0010001000101110011011;
		coeff_log1[8] <= 22'b0001111000100110100011;
		coeff_log1[9] <= 22'b0001101011111000100100;
		coeff_log1[10] <= 22'b0001100001100110000000;
		coeff_log1[11] <= 22'b0001011001000110001100;
		coeff_log1[12] <= 22'b0001010001111101100010;
		coeff_log1[13] <= 22'b0001001011111000101000;
		coeff_log1[14] <= 22'b0001000110101001011011;
		coeff_log1[15] <= 22'b0001000010000101100001;
		coeff_log1[16] <= 22'b0000111110000101000010;
		coeff_log1[17] <= 22'b0000111010100001111000;
		coeff_log1[18] <= 22'b0000110111010111010011;
		coeff_log1[19] <= 22'b0000110100100001100001;
		coeff_log1[20] <= 22'b0000110001111101011111;
		coeff_log1[21] <= 22'b0000101111101000101101;
		coeff_log1[22] <= 22'b0000101101100001001011;
		coeff_log1[23] <= 22'b0000101011100101001011;
		coeff_log1[24] <= 22'b0000101001110011010011;
		coeff_log1[25] <= 22'b0000101000001010010110;
		coeff_log1[26] <= 22'b0000100110101001010101;
		coeff_log1[27] <= 22'b0000100101001111011000;
		coeff_log1[28] <= 22'b0000100011111011101111;
		coeff_log1[29] <= 22'b0000100010101101110001;
		coeff_log1[30] <= 22'b0000100001100100111010;
		coeff_log1[31] <= 22'b0000100000100000101011;
		coeff_log1[32] <= 22'b0000011111100000101001;
		coeff_log1[33] <= 22'b0000011110100100011100;
		coeff_log1[34] <= 22'b0000011101101011101110;
		coeff_log1[35] <= 22'b0000011100110110001101;
		coeff_log1[36] <= 22'b0000011100000011100111;
		coeff_log1[37] <= 22'b0000011011010011101110;
		coeff_log1[38] <= 22'b0000011010100110010101;
		coeff_log1[39] <= 22'b0000011001111011001110;
		coeff_log1[40] <= 22'b0000011001010010010000;
		coeff_log1[41] <= 22'b0000011000101011010000;
		coeff_log1[42] <= 22'b0000011000000110000110;
		coeff_log1[43] <= 22'b0000010111100010101001;
		coeff_log1[44] <= 22'b0000010111000000110010;
		coeff_log1[45] <= 22'b0000010110100000011010;
		coeff_log1[46] <= 22'b0000010110000001011011;
		coeff_log1[47] <= 22'b0000010101100011110000;
		coeff_log1[48] <= 22'b0000010101000111010011;
		coeff_log1[49] <= 22'b0000010100101100000000;
		coeff_log1[50] <= 22'b0000010100010001110010;
		coeff_log1[51] <= 22'b0000010011111000100101;
		coeff_log1[52] <= 22'b0000010011100000010110;
		coeff_log1[53] <= 22'b0000010011001001000000;
		coeff_log1[54] <= 22'b0000010010110010100010;
		coeff_log1[55] <= 22'b0000010010011100110111;
		coeff_log1[56] <= 22'b0000010010000111111101;
		coeff_log1[57] <= 22'b0000010001110011110010;
		coeff_log1[58] <= 22'b0000010001100000010011;
		coeff_log1[59] <= 22'b0000010001001101011110;
		coeff_log1[60] <= 22'b0000010000111011010001;
		coeff_log1[61] <= 22'b0000010000101001101001;
		coeff_log1[62] <= 22'b0000010000011000100110;
		coeff_log1[63] <= 22'b0000010000001000000101;
		coeff_log1[64] <= 22'b0000001111111000000101;
		coeff_log1[65] <= 22'b0000001111101000100100;
		coeff_log1[66] <= 22'b0000001111011001100001;
		coeff_log1[67] <= 22'b0000001111001010111011;
		coeff_log1[68] <= 22'b0000001110111100110000;
		coeff_log1[69] <= 22'b0000001110101110111111;
		coeff_log1[70] <= 22'b0000001110100001100111;
		coeff_log1[71] <= 22'b0000001110010100100110;
		coeff_log1[72] <= 22'b0000001110000111111101;
		coeff_log1[73] <= 22'b0000001101111011101010;
		coeff_log1[74] <= 22'b0000001101101111101100;
		coeff_log1[75] <= 22'b0000001101100100000010;
		coeff_log1[76] <= 22'b0000001101011000101100;
		coeff_log1[77] <= 22'b0000001101001101101001;
		coeff_log1[78] <= 22'b0000001101000010110111;
		coeff_log1[79] <= 22'b0000001100111000010111;
		coeff_log1[80] <= 22'b0000001100101110001000;
		coeff_log1[81] <= 22'b0000001100100100001000;
		coeff_log1[82] <= 22'b0000001100011010011001;
		coeff_log1[83] <= 22'b0000001100010000111000;
		coeff_log1[84] <= 22'b0000001100000111100101;
		coeff_log1[85] <= 22'b0000001011111110100001;
		coeff_log1[86] <= 22'b0000001011110101101010;
		coeff_log1[87] <= 22'b0000001011101100111111;
		coeff_log1[88] <= 22'b0000001011100100100010;
		coeff_log1[89] <= 22'b0000001011011100010000;
		coeff_log1[90] <= 22'b0000001011010100001010;
		coeff_log1[91] <= 22'b0000001011001100010000;
		coeff_log1[92] <= 22'b0000001011000100100000;
		coeff_log1[93] <= 22'b0000001010111100111011;
		coeff_log1[94] <= 22'b0000001010110101100001;
		coeff_log1[95] <= 22'b0000001010101110010000;
		coeff_log1[96] <= 22'b0000001010100111001001;
		coeff_log1[97] <= 22'b0000001010100000001011;
		coeff_log1[98] <= 22'b0000001010011001010110;
		coeff_log1[99] <= 22'b0000001010010010101010;
		coeff_log1[100] <= 22'b0000001010001100000111;
		coeff_log1[101] <= 22'b0000001010000101101100;
		coeff_log1[102] <= 22'b0000001001111111011000;
		coeff_log1[103] <= 22'b0000001001111001001101;
		coeff_log1[104] <= 22'b0000001001110011001001;
		coeff_log1[105] <= 22'b0000001001101101001101;
		coeff_log1[106] <= 22'b0000001001100111010111;
		coeff_log1[107] <= 22'b0000001001100001101001;
		coeff_log1[108] <= 22'b0000001001011100000001;
		coeff_log1[109] <= 22'b0000001001010110100000;
		coeff_log1[110] <= 22'b0000001001010001000110;
		coeff_log1[111] <= 22'b0000001001001011110001;
		coeff_log1[112] <= 22'b0000001001000110100011;
		coeff_log1[113] <= 22'b0000001001000001011010;
		coeff_log1[114] <= 22'b0000001000111100011000;
		coeff_log1[115] <= 22'b0000001000110111011011;
		coeff_log1[116] <= 22'b0000001000110010100011;
		coeff_log1[117] <= 22'b0000001000101101110000;
		coeff_log1[118] <= 22'b0000001000101001000011;
		coeff_log1[119] <= 22'b0000001000100100011011;
		coeff_log1[120] <= 22'b0000001000011111111000;
		coeff_log1[121] <= 22'b0000001000011011011001;
		coeff_log1[122] <= 22'b0000001000010110111111;
		coeff_log1[123] <= 22'b0000001000010010101010;
		coeff_log1[124] <= 22'b0000001000001110011001;
		coeff_log1[125] <= 22'b0000001000001010001101;
		coeff_log1[126] <= 22'b0000001000000110000101;
		coeff_log1[127] <= 22'b0000001000000010000001;
		coeff_log1[128] <= 22'b0000000111111110000001;
		coeff_log1[129] <= 22'b0000000111111010000101;
		coeff_log1[130] <= 22'b0000000111110110001100;
		coeff_log1[131] <= 22'b0000000111110010011000;
		coeff_log1[132] <= 22'b0000000111101110100111;
		coeff_log1[133] <= 22'b0000000111101010111010;
		coeff_log1[134] <= 22'b0000000111100111010001;
		coeff_log1[135] <= 22'b0000000111100011101010;
		coeff_log1[136] <= 22'b0000000111100000001000;
		coeff_log1[137] <= 22'b0000000111011100101000;
		coeff_log1[138] <= 22'b0000000111011001001100;
		coeff_log1[139] <= 22'b0000000111010101110011;
		coeff_log1[140] <= 22'b0000000111010010011101;
		coeff_log1[141] <= 22'b0000000111001111001010;
		coeff_log1[142] <= 22'b0000000111001011111010;
		coeff_log1[143] <= 22'b0000000111001000101101;
		coeff_log1[144] <= 22'b0000000111000101100010;
		coeff_log1[145] <= 22'b0000000111000010011011;
		coeff_log1[146] <= 22'b0000000110111111010110;
		coeff_log1[147] <= 22'b0000000110111100010100;
		coeff_log1[148] <= 22'b0000000110111001010101;
		coeff_log1[149] <= 22'b0000000110110110011000;
		coeff_log1[150] <= 22'b0000000110110011011101;
		coeff_log1[151] <= 22'b0000000110110000100101;
		coeff_log1[152] <= 22'b0000000110101101110000;
		coeff_log1[153] <= 22'b0000000110101010111101;
		coeff_log1[154] <= 22'b0000000110101000001100;
		coeff_log1[155] <= 22'b0000000110100101011101;
		coeff_log1[156] <= 22'b0000000110100010110001;
		coeff_log1[157] <= 22'b0000000110100000000111;
		coeff_log1[158] <= 22'b0000000110011101011111;
		coeff_log1[159] <= 22'b0000000110011010111001;
		coeff_log1[160] <= 22'b0000000110011000010101;
		coeff_log1[161] <= 22'b0000000110010101110011;
		coeff_log1[162] <= 22'b0000000110010011010011;
		coeff_log1[163] <= 22'b0000000110010000110101;
		coeff_log1[164] <= 22'b0000000110001110011001;
		coeff_log1[165] <= 22'b0000000110001011111111;
		coeff_log1[166] <= 22'b0000000110001001100111;
		coeff_log1[167] <= 22'b0000000110000111010001;
		coeff_log1[168] <= 22'b0000000110000100111100;
		coeff_log1[169] <= 22'b0000000110000010101001;
		coeff_log1[170] <= 22'b0000000110000000011000;
		coeff_log1[171] <= 22'b0000000101111110001001;
		coeff_log1[172] <= 22'b0000000101111011111011;
		coeff_log1[173] <= 22'b0000000101111001101111;
		coeff_log1[174] <= 22'b0000000101110111100100;
		coeff_log1[175] <= 22'b0000000101110101011011;
		coeff_log1[176] <= 22'b0000000101110011010100;
		coeff_log1[177] <= 22'b0000000101110001001110;
		coeff_log1[178] <= 22'b0000000101101111001010;
		coeff_log1[179] <= 22'b0000000101101101000111;
		coeff_log1[180] <= 22'b0000000101101011000101;
		coeff_log1[181] <= 22'b0000000101101001000101;
		coeff_log1[182] <= 22'b0000000101100111000111;
		coeff_log1[183] <= 22'b0000000101100101001001;
		coeff_log1[184] <= 22'b0000000101100011001101;
		coeff_log1[185] <= 22'b0000000101100001010011;
		coeff_log1[186] <= 22'b0000000101011111011010;
		coeff_log1[187] <= 22'b0000000101011101100010;
		coeff_log1[188] <= 22'b0000000101011011101011;
		coeff_log1[189] <= 22'b0000000101011001110110;
		coeff_log1[190] <= 22'b0000000101011000000001;
		coeff_log1[191] <= 22'b0000000101010110001110;
		coeff_log1[192] <= 22'b0000000101010100011101;
		coeff_log1[193] <= 22'b0000000101010010101100;
		coeff_log1[194] <= 22'b0000000101010000111101;
		coeff_log1[195] <= 22'b0000000101001111001110;
		coeff_log1[196] <= 22'b0000000101001101100001;
		coeff_log1[197] <= 22'b0000000101001011110101;
		coeff_log1[198] <= 22'b0000000101001010001010;
		coeff_log1[199] <= 22'b0000000101001000100000;
		coeff_log1[200] <= 22'b0000000101000110110111;
		coeff_log1[201] <= 22'b0000000101000101001111;
		coeff_log1[202] <= 22'b0000000101000011101001;
		coeff_log1[203] <= 22'b0000000101000010000011;
		coeff_log1[204] <= 22'b0000000101000000011110;
		coeff_log1[205] <= 22'b0000000100111110111010;
		coeff_log1[206] <= 22'b0000000100111101010111;
		coeff_log1[207] <= 22'b0000000100111011110110;
		coeff_log1[208] <= 22'b0000000100111010010101;
		coeff_log1[209] <= 22'b0000000100111000110101;
		coeff_log1[210] <= 22'b0000000100110111010101;
		coeff_log1[211] <= 22'b0000000100110101110111;
		coeff_log1[212] <= 22'b0000000100110100011010;
		coeff_log1[213] <= 22'b0000000100110010111101;
		coeff_log1[214] <= 22'b0000000100110001100010;
		coeff_log1[215] <= 22'b0000000100110000000111;
		coeff_log1[216] <= 22'b0000000100101110101101;
		coeff_log1[217] <= 22'b0000000100101101010100;
		coeff_log1[218] <= 22'b0000000100101011111100;
		coeff_log1[219] <= 22'b0000000100101010100100;
		coeff_log1[220] <= 22'b0000000100101001001110;
		coeff_log1[221] <= 22'b0000000100100111111000;
		coeff_log1[222] <= 22'b0000000100100110100011;
		coeff_log1[223] <= 22'b0000000100100101001110;
		coeff_log1[224] <= 22'b0000000100100011111011;
		coeff_log1[225] <= 22'b0000000100100010101000;
		coeff_log1[226] <= 22'b0000000100100001010110;
		coeff_log1[227] <= 22'b0000000100100000000101;
		coeff_log1[228] <= 22'b0000000100011110110100;
		coeff_log1[229] <= 22'b0000000100011101100100;
		coeff_log1[230] <= 22'b0000000100011100010101;
		coeff_log1[231] <= 22'b0000000100011011000110;
		coeff_log1[232] <= 22'b0000000100011001111000;
		coeff_log1[233] <= 22'b0000000100011000101011;
		coeff_log1[234] <= 22'b0000000100010111011110;
		coeff_log1[235] <= 22'b0000000100010110010010;
		coeff_log1[236] <= 22'b0000000100010101000111;
		coeff_log1[237] <= 22'b0000000100010011111100;
		coeff_log1[238] <= 22'b0000000100010010110010;
		coeff_log1[239] <= 22'b0000000100010001101001;
		coeff_log1[240] <= 22'b0000000100010000100000;
		coeff_log1[241] <= 22'b0000000100001111011000;
		coeff_log1[242] <= 22'b0000000100001110010000;
		coeff_log1[243] <= 22'b0000000100001101001001;
		coeff_log1[244] <= 22'b0000000100001100000011;
		coeff_log1[245] <= 22'b0000000100001010111101;
		coeff_log1[246] <= 22'b0000000100001001110111;
		coeff_log1[247] <= 22'b0000000100001000110011;
		coeff_log1[248] <= 22'b0000000100000111101111;
		coeff_log1[249] <= 22'b0000000100000110101011;
		coeff_log1[250] <= 22'b0000000100000101101000;
		coeff_log1[251] <= 22'b0000000100000100100101;
		coeff_log1[252] <= 22'b0000000100000011100011;
		coeff_log1[253] <= 22'b0000000100000010100010;
		coeff_log1[254] <= 22'b0000000100000001100001;
		coeff_log1[255] <= 22'b0000000100000000100000;

		// coeff_log0 table
		coeff_log0[0] <= 13'b1111111111111;
		coeff_log0[1] <= 13'b1101011000001;
		coeff_log0[2] <= 13'b1100010010101;
		coeff_log0[3] <= 13'b1011100110100;
		coeff_log0[4] <= 13'b1011000101111;
		coeff_log0[5] <= 13'b1010101100000;
		coeff_log0[6] <= 13'b1010010110100;
		coeff_log0[7] <= 13'b1010000100001;
		coeff_log0[8] <= 13'b1001110100000;
		coeff_log0[9] <= 13'b1001100101110;
		coeff_log0[10] <= 13'b1001011000111;
		coeff_log0[11] <= 13'b1001001101010;
		coeff_log0[12] <= 13'b1001000010101;
		coeff_log0[13] <= 13'b1000111000110;
		coeff_log0[14] <= 13'b1000101111100;
		coeff_log0[15] <= 13'b1000100111000;
		coeff_log0[16] <= 13'b1000011111000;
		coeff_log0[17] <= 13'b1000010111100;
		coeff_log0[18] <= 13'b1000010000011;
		coeff_log0[19] <= 13'b1000001001101;
		coeff_log0[20] <= 13'b1000000011010;
		coeff_log0[21] <= 13'b0111111101001;
		coeff_log0[22] <= 13'b0111110111010;
		coeff_log0[23] <= 13'b0111110001110;
		coeff_log0[24] <= 13'b0111101100011;
		coeff_log0[25] <= 13'b0111100111010;
		coeff_log0[26] <= 13'b0111100010011;
		coeff_log0[27] <= 13'b0111011101101;
		coeff_log0[28] <= 13'b0111011001000;
		coeff_log0[29] <= 13'b0111010100101;
		coeff_log0[30] <= 13'b0111010000011;
		coeff_log0[31] <= 13'b0111001100010;
		coeff_log0[32] <= 13'b0111001000010;
		coeff_log0[33] <= 13'b0111000100011;
		coeff_log0[34] <= 13'b0111000000100;
		coeff_log0[35] <= 13'b0110111100111;
		coeff_log0[36] <= 13'b0110111001011;
		coeff_log0[37] <= 13'b0110110101111;
		coeff_log0[38] <= 13'b0110110010100;
		coeff_log0[39] <= 13'b0110101111010;
		coeff_log0[40] <= 13'b0110101100000;
		coeff_log0[41] <= 13'b0110101000111;
		coeff_log0[42] <= 13'b0110100101111;
		coeff_log0[43] <= 13'b0110100010111;
		coeff_log0[44] <= 13'b0110100000000;
		coeff_log0[45] <= 13'b0110011101001;
		coeff_log0[46] <= 13'b0110011010011;
		coeff_log0[47] <= 13'b0110010111101;
		coeff_log0[48] <= 13'b0110010101000;
		coeff_log0[49] <= 13'b0110010010011;
		coeff_log0[50] <= 13'b0110001111110;
		coeff_log0[51] <= 13'b0110001101010;
		coeff_log0[52] <= 13'b0110001010110;
		coeff_log0[53] <= 13'b0110001000011;
		coeff_log0[54] <= 13'b0110000110000;
		coeff_log0[55] <= 13'b0110000011110;
		coeff_log0[56] <= 13'b0110000001011;
		coeff_log0[57] <= 13'b0101111111001;
		coeff_log0[58] <= 13'b0101111101000;
		coeff_log0[59] <= 13'b0101111010110;
		coeff_log0[60] <= 13'b0101111000101;
		coeff_log0[61] <= 13'b0101110110100;
		coeff_log0[62] <= 13'b0101110100100;
		coeff_log0[63] <= 13'b0101110010100;
		coeff_log0[64] <= 13'b0101110000100;
		coeff_log0[65] <= 13'b0101101110100;
		coeff_log0[66] <= 13'b0101101100100;
		coeff_log0[67] <= 13'b0101101010101;
		coeff_log0[68] <= 13'b0101101000110;
		coeff_log0[69] <= 13'b0101100110111;
		coeff_log0[70] <= 13'b0101100101001;
		coeff_log0[71] <= 13'b0101100011010;
		coeff_log0[72] <= 13'b0101100001100;
		coeff_log0[73] <= 13'b0101011111110;
		coeff_log0[74] <= 13'b0101011110000;
		coeff_log0[75] <= 13'b0101011100010;
		coeff_log0[76] <= 13'b0101011010101;
		coeff_log0[77] <= 13'b0101011001000;
		coeff_log0[78] <= 13'b0101010111010;
		coeff_log0[79] <= 13'b0101010101110;
		coeff_log0[80] <= 13'b0101010100001;
		coeff_log0[81] <= 13'b0101010010100;
		coeff_log0[82] <= 13'b0101010001000;
		coeff_log0[83] <= 13'b0101001111011;
		coeff_log0[84] <= 13'b0101001101111;
		coeff_log0[85] <= 13'b0101001100011;
		coeff_log0[86] <= 13'b0101001010111;
		coeff_log0[87] <= 13'b0101001001011;
		coeff_log0[88] <= 13'b0101001000000;
		coeff_log0[89] <= 13'b0101000110100;
		coeff_log0[90] <= 13'b0101000101001;
		coeff_log0[91] <= 13'b0101000011110;
		coeff_log0[92] <= 13'b0101000010010;
		coeff_log0[93] <= 13'b0101000000111;
		coeff_log0[94] <= 13'b0100111111101;
		coeff_log0[95] <= 13'b0100111110010;
		coeff_log0[96] <= 13'b0100111100111;
		coeff_log0[97] <= 13'b0100111011101;
		coeff_log0[98] <= 13'b0100111010010;
		coeff_log0[99] <= 13'b0100111001000;
		coeff_log0[100] <= 13'b0100110111101;
		coeff_log0[101] <= 13'b0100110110011;
		coeff_log0[102] <= 13'b0100110101001;
		coeff_log0[103] <= 13'b0100110011111;
		coeff_log0[104] <= 13'b0100110010110;
		coeff_log0[105] <= 13'b0100110001100;
		coeff_log0[106] <= 13'b0100110000010;
		coeff_log0[107] <= 13'b0100101111001;
		coeff_log0[108] <= 13'b0100101101111;
		coeff_log0[109] <= 13'b0100101100110;
		coeff_log0[110] <= 13'b0100101011100;
		coeff_log0[111] <= 13'b0100101010011;
		coeff_log0[112] <= 13'b0100101001010;
		coeff_log0[113] <= 13'b0100101000001;
		coeff_log0[114] <= 13'b0100100111000;
		coeff_log0[115] <= 13'b0100100101111;
		coeff_log0[116] <= 13'b0100100100110;
		coeff_log0[117] <= 13'b0100100011101;
		coeff_log0[118] <= 13'b0100100010101;
		coeff_log0[119] <= 13'b0100100001100;
		coeff_log0[120] <= 13'b0100100000100;
		coeff_log0[121] <= 13'b0100011111011;
		coeff_log0[122] <= 13'b0100011110011;
		coeff_log0[123] <= 13'b0100011101010;
		coeff_log0[124] <= 13'b0100011100010;
		coeff_log0[125] <= 13'b0100011011010;
		coeff_log0[126] <= 13'b0100011010010;
		coeff_log0[127] <= 13'b0100011001010;
		coeff_log0[128] <= 13'b0100011000010;
		coeff_log0[129] <= 13'b0100010111010;
		coeff_log0[130] <= 13'b0100010110010;
		coeff_log0[131] <= 13'b0100010101010;
		coeff_log0[132] <= 13'b0100010100010;
		coeff_log0[133] <= 13'b0100010011011;
		coeff_log0[134] <= 13'b0100010010011;
		coeff_log0[135] <= 13'b0100010001011;
		coeff_log0[136] <= 13'b0100010000100;
		coeff_log0[137] <= 13'b0100001111100;
		coeff_log0[138] <= 13'b0100001110101;
		coeff_log0[139] <= 13'b0100001101110;
		coeff_log0[140] <= 13'b0100001100110;
		coeff_log0[141] <= 13'b0100001011111;
		coeff_log0[142] <= 13'b0100001011000;
		coeff_log0[143] <= 13'b0100001010001;
		coeff_log0[144] <= 13'b0100001001010;
		coeff_log0[145] <= 13'b0100001000011;
		coeff_log0[146] <= 13'b0100000111100;
		coeff_log0[147] <= 13'b0100000110101;
		coeff_log0[148] <= 13'b0100000101110;
		coeff_log0[149] <= 13'b0100000100111;
		coeff_log0[150] <= 13'b0100000100000;
		coeff_log0[151] <= 13'b0100000011001;
		coeff_log0[152] <= 13'b0100000010010;
		coeff_log0[153] <= 13'b0100000001100;
		coeff_log0[154] <= 13'b0100000000101;
		coeff_log0[155] <= 13'b0011111111111;
		coeff_log0[156] <= 13'b0011111111000;
		coeff_log0[157] <= 13'b0011111110001;
		coeff_log0[158] <= 13'b0011111101011;
		coeff_log0[159] <= 13'b0011111100100;
		coeff_log0[160] <= 13'b0011111011110;
		coeff_log0[161] <= 13'b0011111011000;
		coeff_log0[162] <= 13'b0011111010001;
		coeff_log0[163] <= 13'b0011111001011;
		coeff_log0[164] <= 13'b0011111000101;
		coeff_log0[165] <= 13'b0011110111111;
		coeff_log0[166] <= 13'b0011110111001;
		coeff_log0[167] <= 13'b0011110110010;
		coeff_log0[168] <= 13'b0011110101100;
		coeff_log0[169] <= 13'b0011110100110;
		coeff_log0[170] <= 13'b0011110100000;
		coeff_log0[171] <= 13'b0011110011010;
		coeff_log0[172] <= 13'b0011110010100;
		coeff_log0[173] <= 13'b0011110001110;
		coeff_log0[174] <= 13'b0011110001000;
		coeff_log0[175] <= 13'b0011110000011;
		coeff_log0[176] <= 13'b0011101111101;
		coeff_log0[177] <= 13'b0011101110111;
		coeff_log0[178] <= 13'b0011101110001;
		coeff_log0[179] <= 13'b0011101101100;
		coeff_log0[180] <= 13'b0011101100110;
		coeff_log0[181] <= 13'b0011101100000;
		coeff_log0[182] <= 13'b0011101011011;
		coeff_log0[183] <= 13'b0011101010101;
		coeff_log0[184] <= 13'b0011101001111;
		coeff_log0[185] <= 13'b0011101001010;
		coeff_log0[186] <= 13'b0011101000100;
		coeff_log0[187] <= 13'b0011100111111;
		coeff_log0[188] <= 13'b0011100111001;
		coeff_log0[189] <= 13'b0011100110100;
		coeff_log0[190] <= 13'b0011100101111;
		coeff_log0[191] <= 13'b0011100101001;
		coeff_log0[192] <= 13'b0011100100100;
		coeff_log0[193] <= 13'b0011100011111;
		coeff_log0[194] <= 13'b0011100011001;
		coeff_log0[195] <= 13'b0011100010100;
		coeff_log0[196] <= 13'b0011100001111;
		coeff_log0[197] <= 13'b0011100001010;
		coeff_log0[198] <= 13'b0011100000100;
		coeff_log0[199] <= 13'b0011011111111;
		coeff_log0[200] <= 13'b0011011111010;
		coeff_log0[201] <= 13'b0011011110101;
		coeff_log0[202] <= 13'b0011011110000;
		coeff_log0[203] <= 13'b0011011101011;
		coeff_log0[204] <= 13'b0011011100110;
		coeff_log0[205] <= 13'b0011011100001;
		coeff_log0[206] <= 13'b0011011011100;
		coeff_log0[207] <= 13'b0011011010111;
		coeff_log0[208] <= 13'b0011011010010;
		coeff_log0[209] <= 13'b0011011001101;
		coeff_log0[210] <= 13'b0011011001000;
		coeff_log0[211] <= 13'b0011011000100;
		coeff_log0[212] <= 13'b0011010111111;
		coeff_log0[213] <= 13'b0011010111010;
		coeff_log0[214] <= 13'b0011010110101;
		coeff_log0[215] <= 13'b0011010110000;
		coeff_log0[216] <= 13'b0011010101100;
		coeff_log0[217] <= 13'b0011010100111;
		coeff_log0[218] <= 13'b0011010100010;
		coeff_log0[219] <= 13'b0011010011110;
		coeff_log0[220] <= 13'b0011010011001;
		coeff_log0[221] <= 13'b0011010010100;
		coeff_log0[222] <= 13'b0011010010000;
		coeff_log0[223] <= 13'b0011010001011;
		coeff_log0[224] <= 13'b0011010000110;
		coeff_log0[225] <= 13'b0011010000010;
		coeff_log0[226] <= 13'b0011001111101;
		coeff_log0[227] <= 13'b0011001111001;
		coeff_log0[228] <= 13'b0011001110100;
		coeff_log0[229] <= 13'b0011001110000;
		coeff_log0[230] <= 13'b0011001101011;
		coeff_log0[231] <= 13'b0011001100111;
		coeff_log0[232] <= 13'b0011001100011;
		coeff_log0[233] <= 13'b0011001011110;
		coeff_log0[234] <= 13'b0011001011010;
		coeff_log0[235] <= 13'b0011001010101;
		coeff_log0[236] <= 13'b0011001010001;
		coeff_log0[237] <= 13'b0011001001101;
		coeff_log0[238] <= 13'b0011001001001;
		coeff_log0[239] <= 13'b0011001000100;
		coeff_log0[240] <= 13'b0011001000000;
		coeff_log0[241] <= 13'b0011000111100;
		coeff_log0[242] <= 13'b0011000110111;
		coeff_log0[243] <= 13'b0011000110011;
		coeff_log0[244] <= 13'b0011000101111;
		coeff_log0[245] <= 13'b0011000101011;
		coeff_log0[246] <= 13'b0011000100111;
		coeff_log0[247] <= 13'b0011000100011;
		coeff_log0[248] <= 13'b0011000011110;
		coeff_log0[249] <= 13'b0011000011010;
		coeff_log0[250] <= 13'b0011000010110;
		coeff_log0[251] <= 13'b0011000010010;
		coeff_log0[252] <= 13'b0011000001110;
		coeff_log0[253] <= 13'b0011000001010;
		coeff_log0[254] <= 13'b0011000000110;
		coeff_log0[255] <= 13'b0011000000010;

	end
end
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module Poly_sqrt(clock, reset, Datain, DataOut);
input clock;
input reset;
input [30:0] Datain;
output reg [16:0] DataOut;

//initialization of registers
reg [42:0] numb1;
reg [19:0] numb2;
reg [13:0] Fraction_bit;
reg [3:0] Integer_bit;
reg [11:0] sqrt_coeff1[64];
reg [19:0] sqrt_coeff0[64];

always @(posedge clock)
begin
	if(!reset)
	begin

		numb1 = Datain * sqrt_coeff1[Datain[30:25]];
		numb2 = sqrt_coeff0[Datain[30:25]];

		Fraction_bit = numb1[35:23] + numb2[16:4];
		Integer_bit =  numb1[39:36] + numb2[19:17] + Fraction_bit[13];
		DataOut[12:0] <=  Fraction_bit[12:0];
		DataOut[16:13] <= Integer_bit[3:0];

	end

	else begin

	//Coefficient 1 Table by poly method from matlab

		sqrt_coeff1[0] <= 12'b100100010001;
		sqrt_coeff1[1] <= 12'b010010101001;
		sqrt_coeff1[2] <= 12'b001110010111;
		sqrt_coeff1[3] <= 12'b001100000111;
		sqrt_coeff1[4] <= 12'b001010101011;
		sqrt_coeff1[5] <= 12'b001001101010;
		sqrt_coeff1[6] <= 12'b001000111000;
		sqrt_coeff1[7] <= 12'b001000010001;
		sqrt_coeff1[8] <= 12'b000111110001;
		sqrt_coeff1[9] <= 12'b000111010110;
		sqrt_coeff1[10] <= 12'b000110111111;
		sqrt_coeff1[11] <= 12'b000110101011;
		sqrt_coeff1[12] <= 12'b000110011010;
		sqrt_coeff1[13] <= 12'b000110001010;
		sqrt_coeff1[14] <= 12'b000101111100;
		sqrt_coeff1[15] <= 12'b000101110000;
		sqrt_coeff1[16] <= 12'b000101100101;
		sqrt_coeff1[17] <= 12'b000101011010;
		sqrt_coeff1[18] <= 12'b000101010001;
		sqrt_coeff1[19] <= 12'b000101001000;
		sqrt_coeff1[20] <= 12'b000101000000;
		sqrt_coeff1[21] <= 12'b000100111000;
		sqrt_coeff1[22] <= 12'b000100110001;
		sqrt_coeff1[23] <= 12'b000100101011;
		sqrt_coeff1[24] <= 12'b000100100101;
		sqrt_coeff1[25] <= 12'b000100011111;
		sqrt_coeff1[26] <= 12'b000100011001;
		sqrt_coeff1[27] <= 12'b000100010100;
		sqrt_coeff1[28] <= 12'b000100001111;
		sqrt_coeff1[29] <= 12'b000100001011;
		sqrt_coeff1[30] <= 12'b000100000110;
		sqrt_coeff1[31] <= 12'b000100000010;
		sqrt_coeff1[32] <= 12'b000011111110;
		sqrt_coeff1[33] <= 12'b000011111010;
		sqrt_coeff1[34] <= 12'b000011110111;
		sqrt_coeff1[35] <= 12'b000011110011;
		sqrt_coeff1[36] <= 12'b000011110000;
		sqrt_coeff1[37] <= 12'b000011101100;
		sqrt_coeff1[38] <= 12'b000011101001;
		sqrt_coeff1[39] <= 12'b000011100110;
		sqrt_coeff1[40] <= 12'b000011100100;
		sqrt_coeff1[41] <= 12'b000011100001;
		sqrt_coeff1[42] <= 12'b000011011110;
		sqrt_coeff1[43] <= 12'b000011011100;
		sqrt_coeff1[44] <= 12'b000011011001;
		sqrt_coeff1[45] <= 12'b000011010111;
		sqrt_coeff1[46] <= 12'b000011010100;
		sqrt_coeff1[47] <= 12'b000011010010;
		sqrt_coeff1[48] <= 12'b000011010000;
		sqrt_coeff1[49] <= 12'b000011001110;
		sqrt_coeff1[50] <= 12'b000011001100;
		sqrt_coeff1[51] <= 12'b000011001010;
		sqrt_coeff1[52] <= 12'b000011001000;
		sqrt_coeff1[53] <= 12'b000011000110;
		sqrt_coeff1[54] <= 12'b000011000100;
		sqrt_coeff1[55] <= 12'b000011000010;
		sqrt_coeff1[56] <= 12'b000011000001;
		sqrt_coeff1[57] <= 12'b000010111111;
		sqrt_coeff1[58] <= 12'b000010111101;
		sqrt_coeff1[59] <= 12'b000010111100;
		sqrt_coeff1[60] <= 12'b000010111010;
		sqrt_coeff1[61] <= 12'b000010111001;
		sqrt_coeff1[62] <= 12'b000010110111;
		sqrt_coeff1[63] <= 12'b000010110110;

	//Coefficient0 Table

		sqrt_coeff0[0] <= 20'b00001100000001100001;
		sqrt_coeff0[1] <= 20'b00011011001101011001;
		sqrt_coeff0[2] <= 20'b00100011100011000010;
		sqrt_coeff0[3] <= 20'b00101010001100011011;
		sqrt_coeff0[4] <= 20'b00101111111001111101;
		sqrt_coeff0[5] <= 20'b00110100111111110000;
		sqrt_coeff0[6] <= 20'b00111001101000100111;
		sqrt_coeff0[7] <= 20'b00111101111011001000;
		sqrt_coeff0[8] <= 20'b01000001111011101111;
		sqrt_coeff0[9] <= 20'b01000101101101100011;
		sqrt_coeff0[10] <= 20'b01001001010010110111;
		sqrt_coeff0[11] <= 20'b01001100101101011101;
		sqrt_coeff0[12] <= 20'b01001111111110101101;
		sqrt_coeff0[13] <= 20'b01010011000111101101;
		sqrt_coeff0[14] <= 20'b01010110001001010111;
		sqrt_coeff0[15] <= 20'b01011001000100011101;
		sqrt_coeff0[16] <= 20'b01011011111001100101;
		sqrt_coeff0[17] <= 20'b01011110101001010010;
		sqrt_coeff0[18] <= 20'b01100001010100000010;
		sqrt_coeff0[19] <= 20'b01100011111010001101;
		sqrt_coeff0[20] <= 20'b01100110011100001011;
		sqrt_coeff0[21] <= 20'b01101000111010001111;
		sqrt_coeff0[22] <= 20'b01101011010100101010;
		sqrt_coeff0[23] <= 20'b01101101101011101100;
		sqrt_coeff0[24] <= 20'b01101111111111100010;
		sqrt_coeff0[25] <= 20'b01110010010000011000;
		sqrt_coeff0[26] <= 20'b01110100011110011010;
		sqrt_coeff0[27] <= 20'b01110110101001110010;
		sqrt_coeff0[28] <= 20'b01111000110010101010;
		sqrt_coeff0[29] <= 20'b01111010111001001001;
		sqrt_coeff0[30] <= 20'b01111100111101010111;
		sqrt_coeff0[31] <= 20'b01111110111111011011;
		sqrt_coeff0[32] <= 20'b10000000111111011100;
		sqrt_coeff0[33] <= 20'b10000010111101100000;
		sqrt_coeff0[34] <= 20'b10000100111001101101;
		sqrt_coeff0[35] <= 20'b10000110110100000111;
		sqrt_coeff0[36] <= 20'b10001000101100110011;
		sqrt_coeff0[37] <= 20'b10001010100011110110;
		sqrt_coeff0[38] <= 20'b10001100011001010101;
		sqrt_coeff0[39] <= 20'b10001110001101010010;
		sqrt_coeff0[40] <= 20'b10001111111111110010;
		sqrt_coeff0[41] <= 20'b10010001110000111000;
		sqrt_coeff0[42] <= 20'b10010011100000100111;
		sqrt_coeff0[43] <= 20'b10010101001111000010;
		sqrt_coeff0[44] <= 20'b10010110111100001101;
		sqrt_coeff0[45] <= 20'b10011000101000001010;
		sqrt_coeff0[46] <= 20'b10011010010010111011;
		sqrt_coeff0[47] <= 20'b10011011111100100011;
		sqrt_coeff0[48] <= 20'b10011101100101000100;
		sqrt_coeff0[49] <= 20'b10011111001100100000;
		sqrt_coeff0[50] <= 20'b10100000110010111010;
		sqrt_coeff0[51] <= 20'b10100010011000010100;
		sqrt_coeff0[52] <= 20'b10100011111100101110;
		sqrt_coeff0[53] <= 20'b10100101100000001100;
		sqrt_coeff0[54] <= 20'b10100111000010101111;
		sqrt_coeff0[55] <= 20'b10101000100100011000;
		sqrt_coeff0[56] <= 20'b10101010000101001001;
		sqrt_coeff0[57] <= 20'b10101011100101000011;
		sqrt_coeff0[58] <= 20'b10101101000100001000;
		sqrt_coeff0[59] <= 20'b10101110100010011001;
		sqrt_coeff0[60] <= 20'b10101111111111111000;
		sqrt_coeff0[61] <= 20'b10110001011100100110;
		sqrt_coeff0[62] <= 20'b10110010111000100011;
		sqrt_coeff0[63] <= 20'b10110100010011110010;

	end
end
endmodule



	
	
